	prg prg_inst(
		.clk,
		.rst,
		.v2,
		.start,
		.W,
		.pw,
		.prg_to_shader_stall,
		.prg_to_shader_valid,
		.prg_to_shader_data
	);

	scene_int scene_int_inst(
		.clk,
		.rst,
		.v2,
		.sceneAABB,
		.rst, 
		.sint_to_tarb_stall 
	);

	arbitor arbitor_inst(
		.clk,
		.rst,
		.rst,
		.valid_us,
		.stall_us,
		.data_us,
		.valid_ds,
		.stall_ds,
		.data_ds
	);

	trav_unit trav_unit_inst(
		.clk,
		.rst,
		.rst,
		.tcache_to_trav_valid,
		.tcache_to_trav_data,
		.tcache_to_trav_stall,
		.trav_to_rs_valid,
		.trav_to_rs_data,
		.trav_to_rs_stall,
		.rs_to_trav_valid,
		.rs_to_trav_data,
		.rs_to_trav_stall,
		.trav_to_ss_valid,
		.trav_to_ss_data,
		.trav_to_ss_stall,
		.trav_to_tarb_valid,
		.trav_to_tarb_data,
		.trav_to_tarb_stall,
		.trav_to_larb_valid,
		.trav_to_larb_data,
		.trav_to_larb_stall,
		.trav_to_list_valid,
		.trav_to_list_data,
		.trav_to_list_stall
	);

	shortstack_unit shortstack_unit_inst(
		.clk,
		.rst,
		.rst,
		.trav0_to_ss_valid,
		.trav0_to_ss_data,
		.trav0_to_ss_stall,
		.trav1_to_ss_valid,
		.trav1_to_ss_data,
		.trav1_to_ss_stall,
		.sint_to_ss_valid,
		.sint_to_ss_data,
		.sint_to_ss_stall,
		.list_to_ss_valid,
		.list_to_ss_data,
		.list_to_ss_stall,
		.ss_to_shader_valid,
		.ss_to_shader_data,
		.ss_to_shader_stall,
		.ss_to_tarb_valid0,
		.ss_to_tarb_data0,
		.ss_to_tarb_stall0,
		.ss_to_tarb_valid1,
		.ss_to_tarb_data1,
		.ss_to_tarb_stall1
	);

	raystore raystore_inst(
		.clk,
		.rst,
		.trav0_to_rs_data,
		.trav0_to_rs_valid,
		.trav0_to_rs_stall,
		.trav1_to_rs_data,
		.trav1_to_rs_valid,
		.trav1_to_rs_stall,
		.icache_to_rs_data,
		.icache_to_rs_valid,
		.icache_to_rs_stall,
		.list_to_rs_data,
		.list_to_rs_valid,
		.list_to_rs_stall,
		.rs_to_trav0_data,
		.rs_to_trav0_valid,
		.rs_to_trav0_stall,
		.rs_to_trav1_data,
		.rs_to_trav1_valid,
		.rs_to_trav1_stall,
		.rs_to_int_data,
		.rs_to_int_valid,
		.rs_to_int_stall,
		.rs_to_pcalc_data,
		.rs_to_pcalc_valid,
		.rs_to_pcalc_stall,
		.raystore_we,
		.raystore_write_addr,
		.raystore_write_data,
		.rst
		.us_valid,
		.us_stall,
		.pipe_stall,
		.pipe_valid,
		.data_sel,
		.mux_sel0,
		.mux_sel1,
		.raystore_we,
		.rrp
	);

	int_unit int_unit_inst(
		.clk,
		.rst,
		.rst,
		.rs_to_int_valid,
		.rs_to_int_data,
		.rs_to_int_stall,
		.int_to_list_valid,
		.int_to_list_data,
		.int_to_list_stall,
		.int_to_larb_valid,
		.int_to_larb_data,
		.int_to_larb_stall
	);

	list_unit list_unit_inst(
		.clk,
		.rst,
		.rst,
		.trav0_to_list_valid,
		.trav0_to_list_data,
		.trav0_to_list_stall,
		.trav1_to_list_valid,
		.trav1_to_list_data,
		.trav1_to_list_stall,
		.int_to_list_valid,
		.int_to_list_data,
		.int_to_list_stall,
		.list_to_ss_valid,
		.list_to_ss_data,
		.list_to_ss_stall,
		.list_to_rs_valid,
		.list_to_rs_data,
		.list_to_rs_stall
		.intersection 
		.logic
	);

	scene_int scene_int_inst(
		.clk,
		.rst,
		.v2,
		.sceneAABB,
		.rst, 
		.shader_to_sint_valid,
		.shader_to_sint_data,
		.shader_to_sint_stall,
		.sint_to_shader_valid,
		.sint_to_shader_data,
		.sint_to_shader_stall,
		.sint_to_ss_valid,
		.sint_to_ss_data,
		.sint_to_ss_stall,
		.sint_to_tarb_valid,
		.sint_to_tarb_data,
		.sint_to_tarb_stall 
	);

	simple_shader_unit simple_shader_unit_inst(
		.clk,
		.rst,
		.rst,
		.prg_to_shader_valid,
		.prg_to_shader_data,
		.prg_to_shader_stall,
		.pcalc_to_shader_valid,
		.pcalc_to_shader_data,
		.pcalc_to_shader_stall,
		.int_to_shader_valid,
		.int_to_shader_data,
		.int_to_shader_stall,
		.sint_to_shader_valid,
		.sint_to_shader_data,
		.sint_to_shader_stall,
		.ss_to_shader_valid,
		.ss_to_shader_data,
		.ss_to_shader_stall,
		.pb_we,
		.pb_full,
		.pb_data_out,
		.shader_to_sint_valid,
		.shader_to_sint_data,
		.shader_to_sint_stall,
		.raystore_we,
		.raystore_write_addr,
		.raystore_write_data
		.buffer
	);

