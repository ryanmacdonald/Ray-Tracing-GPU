module intersection_unit(
  input clk,
  input rst,
  
  input LNT_to_INT int_in,
  input
  output INT_to_LNT int_out,


)

