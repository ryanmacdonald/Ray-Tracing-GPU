
module BM(


  );





endmodule

