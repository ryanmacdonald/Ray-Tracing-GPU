// OBVIOUSLY THIS FILE IS NOT NEAR COMPLETE
/*
module color_convert(
	input logic clk, rst,
	input vector_t color_in,
	input logic v0, v1, v2,
	output logic [7:0] color_out
);

	fp_mult fpm();

	fp_to_int fpti();

	logic less_than_0, greater_than_255;

	assign less_than_0 = int_value < 0;
	assign greater_than_255 = int_value > 255;

	assign color_out = (less_than_0) 

endmodule
*/
