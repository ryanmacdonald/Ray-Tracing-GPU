module trav_math(


  output logic [3:0] trav_case;
  );

   


endmodule
