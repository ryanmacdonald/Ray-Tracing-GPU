module shortstack(


  );


  // Make sure that the entire stack gets cleared when a new ray comes.  And that no rays are using a stack
  // that just had a hit.
