// This is the mailbox wwhich is a memory struture which holds all the hits (and or misses?) that
// occured beyond the leaf node (stores the triID)
// before an intersection is done, this mailbox is checked. If it is valid and find 




module mailbox(


  );






endmodule
