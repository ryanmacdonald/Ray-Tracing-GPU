

module camera_controller(
  input logic 

)
