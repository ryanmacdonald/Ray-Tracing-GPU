typedef packed struct {
  logic sign;
  logic [7:0] exp;
  logic [22:0] man;
} FLOAT;


