// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cfFBSGhPyXMeUznRtXvvBCdsloI0s6CnUdq+ImaOIZv7kbY9BU+kNF1HQjVy+KlE
kV5r5OwP7QDR1KJpJU29eUv3tSNISmzZfoRn8doOaIWMr4QLSrbvnPv9FFK6qjyq
RqyNOvIoNWhZnFA9IuWRHzuN28WLlp961KiVJO6T2UY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 751504)
RqHZAgOsVyl+RCW/MvgfKLZLhSXlfp3XspsJM4EPtjHTBUlz/MBC1LlSI7l22eAO
DQA9GxJdovJ1UHIHJlgXOgZtoSk0M6/tuCWT+UTdfOZdyxIC3LyTzsRmktehv4GR
q1HK+0aPhNKO9cWOdAQkgtnTG59vJ6gZ74fp0P4Vpjvlv1/cdpirDri0dO3hhY4s
a5Ohj31uPEC4Sy2G8arzNhnoTviwiD5phYqQcPv1iMMC3f5K9bIEg80/5pbbO0tK
KPYXitfS4uyi/Nx3iv8H0eo3bF2av1JmJymQqvNM0HPTul9eVnDHKbix7jwwIy/3
05HkCiKm+Gjvd+BHTkEg5mRNzSa//x9b4z8PThpinwLrzUpm4hUcQ61h7owIka8P
iPuEm5FRnyNP1LScdhoOOXmBIxQJacZgK3v1nowR1iGuR0Ow6w2z0bckO9JSCcWG
Lixrzg3uD85RhnY5vJ8Kpq8iJISWitcZdmRMVnEGUzPgVt5iuaum0sUD7ySue53H
ZBdg9CGRnN+flLOmA+GyrJeNiRSJk0pv8Rks7T7s8mtZP4U/yKiesSSXBmI1lisU
ySiJ08zkiHUmu/89FK26rjv7i6jV51YClFeCieI7sonlpMddTozh4QQ/PjCkNs67
+QqPnNad2rp00CQ3CBBkmbfZm7p3+KqtY/kYaiJ3BgfbVfi9xx6DpI+fSwUMiQDL
4u6ZyQDesKcQ+T4S64n6ELCR7FRaV9O59d9wATrrTW1Mvtv71PLeV8U953SWOLxm
F882xQBS0bTJjZrrik3ry3WGsnIFgwXV5bkBtRHz4qAgF11WMKMPxl9oVQxnLmTd
V+V89LmtEDn7nct6dvwKUo3Zmq4IFt2eWN96GzwX9sxBbhW7nv3pwQ0HkJmv1NpP
wcxLmarz8VygNdfuRp3WukSbpPCWMRREXaPh4HT24+FJos0kLeOjwwuca6fKmOOt
KsPEvgrocQlEBwpxcZuxlN9h/+TzLL3IZ/msOaq3FBgExfOig8cifNTCUNUShGrR
HI6LzkygZtEx5pZJIOxNqHxLqjYexI3vucRmuBvlZ8dHOZDkD4SCDhMSaMSMPm1Z
fXAs4TrJRiThB26qZFzGpHY5+gqEqXwM24x8l5nMZOiSnys2PPIT3gkcNg9gZJlU
yqtm/Ug5gBzDIWDyRZZwYKoqlLZYqnFV2s1oXO53a6XxR4Rae9hNUSPGqWiv2i2g
bX0dFuEZEpsgw5vAx5AXHz+jrDbuyCA0RteFJsBIhJWKNKL3FyOphvVPN4UJ7EC/
5dPCppZKH6SpfCccSU63IQvL+TdfJDve266ke/d2A6ZXq6GOi/FdICs6vNqy9nP3
9nRCtTlW20H9KDrB26wX6SE56GUWk+6S9fipAZbcziLNNij+exiW0LvivK+crvlM
jM5p/hhJuhxlFgO+N+DBaRQO/Fm2Z9NXEU55jt0SvjUsBtqllEwRBSVczPvfEGjb
EU+5j34zbx9n5y4i52PRlYf5nm6MdBcPAkyCjPvEgJrFYPjnyPvc8ejwlWjaIxN0
+FaYJWcH8LfeqpNC1BIgYcSPTDZAs81MNTgPyKO2bYot+DNt9ZlKlEIsXtRe4SS5
lt740Gp3jUXCIcicQGYKfTHIn2KGJwszJENhtOg5lgRQa6c8d/QBcdKu9FbBX1de
Z4QDlAI4bRZckT/Ykkc+Hrns7oTArvdhJ4ihMO/PlWYWJ10leDHmOFp1w5TkJWMk
e+sMZt53aMAh7KCR0yqNFvx9zFN137g3oguR3t9S5hnB9am7eAnBnF9t5oGPbvAd
yoR4/RgvH0RItufqc2ifzIradUY9nutJdfPuZNO4dQ2Bl1pXaudUA1gJO2lDhTF+
lBC5LogTCkEbhZYJZg4girRxl6q/ugKpWYthS/UqGXnc70EXzVXaFT5hUdOaERCh
t6ulGN/iuql4HbdTaNAHbVK/caTnRy32MZV3nz0A2iV1XUupQk38NtAnzcZfR+Mq
WzT/OFYW31SuRTXVDq9NuSlGzyWrJIIE06ySZbV4dIXRZ+xaNxP0iN0dtlyWgQIo
kjfABBlwcKYaW+h6HPBEpHTtlHWfqRuD9lba3c8FWutJmdHI9SGGrrmfD6430hcn
VaPX4AxNN2hzS4tJey2q4KktePGPHTKI0u6YN/vdBCGKk7jwhcYGS0miWS6LkmRN
kYAtL6XxR/ltuFUkw3XyuZEbNlebiGBAJBJD7qc5HajGC/ydJFNfeYX2mzMXUT9H
GfMJVbqdS/TY5Mpuccn/Zxt0Umus7sLp5/Uide1GIOoWJjvYR4gaG4/pNFZGYc/Y
kuWXcmdV/Civ0b+EehsHtc5Uhw9vyVzqAxL8jigjOW752dO1lihbE5RErr8UJmLg
a+kfVCfDVxkGvIm4ytxuiOYwlUtL44+nwsvUgWpEYZYLf+YXxPUQVdbG+/D8q2UQ
7NHvfxAelLbJWiaKmAGM8tOE4XI2qDucph2b1HzhmnjRCafF5jpSDNiusUhGApJv
XeJcYKGAtpoq5v3WNmGifeYstRZ2PthYHaBs50vzbajMAknsf7WW+Cmdu9vyH/BM
cP60NCKnHT/gkVMUNAEL1zmt/vRPK8s3q+uFbIcsJi/PQeHCNZIeoV9RvxfvAAFO
y62EEYFr96BesbIshUknG4dEutO6hq+Ab7iycOBFgrPIlCugHTK2XZpMrMtPUBiE
yijt/UkixM+s/wzIP6ymGC/sfvOWCcdUpsSOlE9xFND5LHZHydtDg4Gf2yOPPJ2q
QW2RH3gBf05phpK99ugEzgJy2DOCQJDldH7It3GAEAYMtL/UXuFPrWM5BbRIB62d
4RVbO5053A8ZE+0nnEnXA9O0idD55/JfIRGy7x65FeukbG9jVIBy//3DMY1AgEx6
zKaZzTvmeL3vcuIuLh+PeEOamVgXq+Gtl3/Cs6XJAc9vinanqJxfg3gNL5n3SJSQ
SpQhSQBFZXX+e0JwpqPvsqE0in08rBiNSYj+1OWmXSXunmUzj6QV518pq+ngxH1X
Q2GY/L574ctMHeXumtgNJHpRCvnuWX09ZmWWe9X5MMH41sHk5b0qAhxMt4R9JyM/
kYO6nWViehzmq7KDkquURC26UgK/ZentatGGs98Vh5oxMeqpOWiK0BB/QeSAKtON
fVEyUdf8T1ZEv1FhVBqYTAoNKxgAvSxza4xtNe+KQd/Ssg+UB8jXur27m7kUc6eo
c7lNxWeMMbcVVdGirSoSVxm2HCLvpH1bv+Q5J4TjdNfcv+Q51W3MKePc8OWcWt6d
EMaL8Spv4htMq8qPec1xEvRV2NOI1w3+tboWihzN5PK1+kX6rKVk5yxSImEHiv4y
kJMYDctFywlccyDY2FL33Wji4vhL9rs272oMt58KW2nL64QZZyoV9xRJn5/sYcUh
JFvxBGKCFy2hbit7f3HS2YVZDoHjyDw8M8zwnvs/7yyY1IfVDvaT7tmBF1CkNL9p
jaPdMF+UW0ewu++LCplvj8oWZEz1+oPNfV9lBJH55/YhLQQmOpaU1mKMZBUz8cPW
0fSXnPSZMv49iYS32KZgV/n43oX4pl1ydiEvODp8i+qN+wAU2aCAmRMWDOcSCXaq
2a4z4dbPN+efmmxVnXlulh5N7G+zQDxnPzP0bbAhobvc/ba1doFsJcsP2W3Kbc/s
GQ5zmw8e4nSMLm/hMDVrOXkM7LG8WDk84MvzknyP5HDo/Pds8cUvtFTdPpj8gPWV
oiEZBe44X0H6zoJM9LBANQXaHtMuq6dQGITkA5lQESZw3wtQgiSMgp9BU66oKR3i
NJqSMYMoPxXGucLG25jdfWyJn3POB16g5Xxhroh56HisxybMKxaZYeft8LKEHDzs
LsMa+l/E2u/uOEq0hoeSZkhZIQRCjlti4CgAWlp9vIc5510xY8u4nvrcTzYlTIVH
MpDlBz+1bg0VRwW+TD2ORcvFowotAFTMt+abJVHwcJQXWVIXo4X4y7E2E2KgZfA4
e2+Z2O8oJV6LBtVuRxiFcmcP3yIpDgNq3CZTwmUxVWeBAgDwg9upFBoSrRmzKQbo
nyfIIw3qNefvZ09XmYqAAdu7udNJL8ccXLX3ox8t3rxNKQg6zFOROGS56p8zd3bZ
7bAg+bGUxXpMW5NmjKsceo3dmc0SDUdnGWBFMhc2xx2Pt+tMfD5id8q3HqsWmiUW
5yR5XIQzd3ieh5vMeKlDZmtJn2NrOYqW9/fjtZ23M14qxWOD81/4U34V19wrpIHA
oje/hcS1x20Gy1GtKenLvMfn9q//r+N+3qGZl+7CQnWHOcd3sKBBkrnQve2fYBSK
QM428LsinTzCl0R6/iQgqAJ7DzfJAaemD74M/AUGeyV7gqwBVj0PnXTJxbQkr1ig
J4Ub8AnffnfYoyV1/BuGmIZ8u2Dg7Ax0bF9lRvQML79EiXB0ZHJrkMuEQ9LtwBK8
FJpOowXqgf49JgFAPqiLaPabqzaU6BvTfjWATA9rxgM9KmiYnhJfK6VQK3s7YO2d
AwpIUJLotz/X36bZnTzctO8TzR4bZlHK1jl7huB/rH1bVespEM6hQYslYcWnhKoA
CntUK8yxJhm2TyIsYM+YqATVueuBhdFzzl3v7x7OOOo4hShi7yOikNDDYE4OKrJ5
YAb9umf7oHEjQoluAg29P3q9jnFYjSpLmv8pCfwulZ8deGd6fQeiW428c+io89p0
Q95XLplesoxEVTcrEhXt3BAUjDfb0N2uCkqWMmO7mzfSXonF8AyS244k5IDPvW20
vHrO4TTtB+trSbQaFk+U/mj2axfMFoVr3MieXopgyl3DUY4NY/QS9RWTdXv9LSLZ
KMY5ecqLIqfu589yU1fiEBZN1hsgfBF5VzohQsv5AqaTqbQvnm1xdoSu4xIiZhxo
hH1MPo7kVzeW2hXxv9lhuNt4RPePckG9NaW+SPDDtuWCfRhn7YNn+wF3MBLCmIWb
f9UPWmoIrGFwyUXjyrVsiJttXYSZ2BGDaKPvvOCRwvgfw9UTNEmhpa+t8E7s1hSk
5ocijItXFPNe13oMQheDnFPKuKG547thrcTwjRb3P2qI75ogW9+z0mbhfdApgi3E
u8F0JI8ivcLNvjPhuYq1tSOx8pbYvhnQcRXYrgJDA/dyoEIn6IZXqozsQ6LfcwxN
++SzEH3K+J/eUUGI9b+8dk7cOBpD3G+m4uE6LVwnvHz/xUQYjKiGH3X7/g3kZFFa
7ZYjmjAIH01YlinrUzd82R10uQU832mz+nln0yCQEDXssjzEOBa2MZ58BXYPuwmL
Qm12dmHjZV730mr2NWAHAFLL3NxWaH+Y6XYLgEZGyRjPgwns5Wc+51JQz2xBJwFc
APAjqvqOl7JVofburqbHcsZrEmGqHMVBXhkjPAl1On5YqTInKQxM6YRqZhZXuoBH
WdmJjTbR35lfVj0rMdFARiQAPi74oqHc/byO8RKRfYxFAAhKIS6eqWXHko9HdNL1
b7lrHJlnWBs2Z91QM8/3Gy70PijN9BJjrYXcLIO9SRjDCesRPyq21aS8PPlPxIC5
Yh7EGbaFcEbFVFYbGdNbP09JXIz6QgM/YAe4D6M38L6uu3w+Qo2VY6qHctsHQw93
13TXApLRC8sfQULm51icRz0+G8+Re1LlTsQQqLjhbBNc9abLJJBWomuTTwoK3hcd
Um17Yh/HqHmHioDM6dmx9IP6lziRSCUqAi2rPDoQoRYQ9rf0BMELnwzObR1VTafI
XqCwM1hH6STJriUizXSr1XhVrCmDq/V/Z2ywkGpZDk4LTlztacQu9hh8Kxpf1BO7
PX+6E7MB8av8442YLqY1UqrYPNmXTuIez0UYZ3qJKohic+fXx7bFZnd0rbKXh28N
RzBWETYnB9V6xwM5zGW8XQyGUo/TzhndurHdZUtJWWbR9JGXLNGH3S5Pss8BKAYP
3fUJUSKZ7yfKVBq5x3OhWwhmnqiNvPLyhFc1Z1rlAgZZasIl0iCmc2xVubD9XuZ5
AKeRa17cPo9Jgmpbsq4/DUUIQXWX71wzUnnaiwSnq987O9qPEjq0Qt3GxeXw83d+
/EUL5oeA4S/MThnWil+hSeOhpaOnsDiBgI6Ms7CzrlVGhuQo/M38X9QXpTE8wx9F
0T0zCSsdptrPJLWLz1onIlthoYF3rjMRfcTLceEekXH99y1NxZjV5YMy4cbCOaAF
WTKnA4Hi7uBSbbQYd0OfifYdH+Hy1/bDH7SBTfds+lQiAVDtleUatuhQPuHJKCUk
B2LByPohQwAfO0LAeSNsAXPpbDS1GFEqywnn+jB1V9aSlOr/ApxAV1DX3749AS1v
oAqkMBxW4N+TatNNLMM2N9+Y7nZ93ast9tLtpEZQnBIhhFJPu+nh5DH8jf4Kuc/q
LYuZsUDv3J82BP0ctNJ8ncPdXrXA+YBLKZrFbJh9OnvUIZtVaVOntm3r2/xKZM7f
mXFCYKK3JxvlqWE/OT8i++qwyIKLLPWPieA1++e2NRFNxs9VgJ4yFltYjW7osZ3e
8SxNFnCiyE5ECCATXvqVA7D0mbJu5OcruRb7Es7P3UOjg3c53xKnooqXO6GwuHOA
ncxar7YY1OoYA4kU+FilyOuerZvqPvNOM9OK9+Itx9y7QsLg6cyAtjKhEdIUHyjc
/5+YAi2HxY9DP+6gsIIttWc+X85K8GNge6DuDq28Kr/6MQCCgsJ3eP7gsL970/Mr
vUUPWu+ftEAWSxO1ZomsTLR5x6rMDr+QkQJ9FWopnGEaemwNZd1qbEqRGty5AidX
DQ+jNx9WsQA7XkjVCjv+A6QQEwo/7EUKw8S9Z30kzhxA+W7pomOAIFTh+o10cZHa
dBxoaWS+2PvB8ujtCdLR2PFcfnRcvHS6jE3mEKM3dPcTac2zhiLpi2Zb6xSt555C
yNNwQVKtfL02BouFxWwU01/M/J0zX9OJXuvk28+E6YuyFjvbutlsnNmwueg8D7hX
Jx/2r54jZVGxHlUTSHCEqrc/FUfwQhabxYRbR8MNN+0Nj2afBtsq54kGkw/5RbYl
tAP2gM4BlGa3K1Og5hgEuBnYEO9q8ZfD6bu0LwhM490aoNGdSKng9ONOwmPcbbwm
OwbnOeJmephPaiFltLQJjIsQC3GgnZpuIOqnstmik78vT9k9oYsrkLc/lfyZx4V5
e4NJ1IsAbI4ez//Wji+kdrtOifJh1oNHR/+HUkranLXNPHsofz/+KF2dTyJoW7fz
HOJLIkYf4V53PFjyFw96d/rKBZMBv/lP/pjT896EG1bNrm+LW4rivCgx59QN8Qzv
EZMXJ4b3xoG8qJbw7plZAETvwwPC3JKeUu4uVYL5jUWxOOxJyGILz/FikZecSs/b
FCBrAK2r3Y7riqhgWkv0/L1Ad+OxJ/TBbsvhShAMffy7lyTKFtBj57tx6Az7+9wf
tu5TF5t1gtkEXz+3u2qAxlyzGLv71L9XJ0kKdMI8BUk6Z0/FbBKFFonQhN12HvHl
mklH/j6Qj5ej4ZdYb0/yZUkm/jhPKEpArretSjR8vXhWGwfqe1nnf1h/Ukmf3iMo
FKAabpGRQxTOlCXXpUcHCfv1ykeLTt+nO5oR7GOnAPiCeZ6Nlh2T02/GV/4ECdjo
wJwH51T3aV2LRDm2SGOiaB7QkDUd3GGJMtZxBn1RhWy6Q1f0ISsHmkWEZvOigpIv
TL8xK56ItzXkcWPacWG5e0exWgCfJnd6MnOV/10tWb151GC1MfmSaX6L4CtNh2v4
kI6AviOqcIeLmqpE+Gd1kXYZR+1mcf6nwJj2C5jxLhtgHZpGKusFgQ6HI3VnC9kG
XhFws4LWEm34uiKlY/S5KZ/b2y6cCriJOk2MMVp7TLnMXlWm/SlPQyP7Y1p7Mr/v
YJYyXMXu9mFAuPT44rDg1GBuCTiKFrVKAu4AodHKH0iR1GIpDnAGyHxzDK8n2FLz
vdq28PzvHiowg/m998/VKPGz9/85LG3lkF3IlsioPCp8pwU5EM04ibo8K1BwCXBJ
tW8LbTkI0c0Zz59sXYwk2WlydsZ/KHOrMlw2kjp5yvB2/wFMx5su3PUrhcbtKMgf
CGLPQ2gpbUwkyOwW2ba5J/parBA/uU8RbgLF+MWNEIAM8tcjh8KL+jqdbD9QZsEm
06iPM7mcIZC3A37zrNlnUvA4hGv+ZbqQ0Mdv5VeLcZHvx2PO9AqrnbrOfuOU98/5
kMuvhtDCWffbig5Rervdnm3RKZa1dLKDY18NF+K6yW2zTbneMJD76mmGq/0VZtY/
SQQJO68zzllE7bVzY0fJ1J0hbk5EwpOVRYizDXqpW5UcPatl/3JlBj8zHis0BEmY
b69p9dEk+NoNlmjFilzxbzvNd2sKlUl7jt/6Q3h+vNkrwMEmGxwXALQMV7hwH3z+
iyFsQ5KQuDz9y9nBvgmi8hLI3rI6Z3xL5oFlH1BxNXYUpGt4PUXKZ41p8DqSYiYz
/eyVWefIAIfCK5uXdUkdhbTX3tfgKPjz7JFbqje54Gq2KivH6P5xd88Ow4bLAqFg
WdP04KD+IGOOvTVP69rFb+KwOnuPQiPXCnukuz8VcFuueqssAfijZ0jgRhHPgQJ0
NtShhh3NMZ+IrkDBVfhe+VEXFwqlYFhmgX/cLI69loGXfaUS5/dWZhigOhNrwkCz
hKhmL7sIv23aX4AStHt145yl+9A9es6E6nMB7pMf3+fPI3aHiWMdhKDLb8RnsbQm
9U+HFk2WF31vKhSffYWuNaX9TJnSVJ4tBcf1N5RQqLRKYH4gCYjc8I9TEbsLWI/a
v85MVD+49pGlgqlxcTpZ0xt6gmGyAEKLzviPFziLgGaTMwy3VL+53xcVzkrwsEEN
byafQCIUYfvBGFa7QopMCU7oZUFt65s6Og/pfsUXXbbQkAOMZWKCXc+uA4fCX3e4
QvWN7EIdKOPXGjRi5/WW+OYm8WpOYxNzExFVoIEh5XPHvmzZCUCHPwKuLDiV8ERF
8HTg0mDz9NqXTexb1mRW3xscazbyPotfiiBYG+pTewuwWNse4/IMrOOMcpfkxoAT
k/SS0oGPf6wj9gJEi/TuqyUmeieia6jf/E7pt6y0La0wn4a08lBPqxYW9zRx/ALc
GVTOTt00GaOoC0LDGB992Ms9oAqN0u09FKsm+8drjuCyRemENpx3WZG2NE6VBp5N
zId8/ZkHO1KDvpihJbamDr0BLU/eRGlz5fY9Xz5vmUwNlK7hOkVbskZg6tl7MOzD
oUPgiYwDsWFm96QJK4tfiWaQv6w+0W5Oqa821BtUKPbUeJpizBl/ByG1YJajh3L3
QR1/2ov5Kj7AeedyKdX3BooKyTqpfkbRrqddocTlazi2oPznt/HKUY7BrzWzyUJd
oSxaqXfEwvv617sa2ci6hhZWxQ4gl1xEalg3DI357Xyt6/5gk9T8zYnoXeVhuCkh
vvV6B+IMgXLmiBgkM8GwFd3c/VEnIrwzII9HQ1XqwC1c13crcJcwrqe4KGT2eaEZ
Nxko/bhYmNKYq3bfeJuHI3Mud0NixyJ5A6/oBRuwJMhRwq8l+jBLVbAAJRf7Y036
mQ5ruPb9mG3Z6gg1HJrrI8xnp9a3tmu8w6ukFQRHtSrIL8BdMvbGE+8e7gDyEG//
/3JI5xnmvTxWa8Sy0RHW0WsB6G9C+Oa+YddyvIBPn38/4EbJ+e5AKF0tr/lizJ7J
VvRLHL6Ql8ijpoeJF4zWx8mLykTR42zj4pV3h33EzqX0Yt1UHw+gHHMICUC05V6J
OC4YbOXbcfmkFBucDP/WabeuBL7FrAfOk+igsQTpji7SyapsgfQA1+IQaHFYycdo
Q89nyOsiqflhyNi5HG/cMjNs5Y03pfb9I5amU4Ne7mtBZn5izyedRkTa1p+TiPpo
wN4VuUwwh2BKghceZzafkcEzXaJclPRmUbgLpt3nxcvhRXMWtY2ydzs4TQy80AEW
VxuWjXbfAQAmj5091D6805vZW7sAesSfEFUrKgJSaI7G+XySfk4PiSJ3j05L+suF
Fg3TS+/wVcoJH6r8GrsywVwn6aJB+K4Rk8P5cyNiwZufdDaKoL0IbX1eO0LPL64m
NOdBAOTSe1nnHAz5cbFWLJA4Ubqqj69UFdnfPXpASfot2oR4KJ51ookw+/n2gNlJ
6vIPMe61y7Mr9zwZe3ywQYSndnY5+V3lBEXQM9xtOjyoGEAJV193QzX3loR5mhIM
rP3Gfk3abwFFc0+phVqCZ2lal6KF3Q1ad7WMwf1VunuHq+PVc0XvcFCfxXJVg1rk
uRotZhpSd3AVCMuFhxBI0854VBIPb1xNbBsX55XKpFq22d5vkABTRwJMhI+qZI+Y
9xmo9c1u862/UowF5LaBE2oT1GjPDYrl7q26milPoFfTZiTAK24DzniGH9tTEcaa
kqZ99molcy0dkxWS3feINF1gLSneJ5/UbA0YMqsvPwsvaTcuSsu243ZZR4iHC7qz
7kGIWE898Ip8+spPIudm0zr6/J55uKFoqabVL5rshskBIx9OxPD8bmiIZCRgvA0m
mP0HFKquNYrZmnWWWJnGBSaP4nOUs+TIx+n4y83M+2RVvbw05fxa1iisd+Q/KziR
geCH7lkCQXwgXUl5mz+fyZj0B2AnLN0eEfEN8oz8FaNlBMbhTBhDpX1ZzRf/hZkI
9pqrWjmWjyS9a0PxUAjSyaeDEfr+SvD6PCOQN2h5SqIPVomYt8Om+PlqtkLwoMPG
oisbEZCrRYbhxPt4k/cU5qZxq+oq6IUv9tXWILU0DjLdSnkTQW5wTC6yeto80P62
OUFLJaaVKgQk2A6yDV9JjFsPvnI36f/9LNUDDADwKOcCnokVp1eT7kVamrfYYD8B
G3jFchuFGvUWxr7agJI5QM484OdyK7dOXs/gVCIFXatJ4tpXmciRle6jhRpP1/ud
jmuDTWMKbA98LTBVLuLEHlrNB9RPY9CQtAOsEo6VfBM1EPRZWQBzQRMZBlnUdfh/
yj0D6/Jm0wmc0c2J6klnznGThXRuRN4YVaRzxVRJA1IlEPpYr2mViwjNUiGeLK5V
2PdLo7u+A0NPvObzgs/aUtg/G2tAz3RM4Doz79gUVefeOkUaYrSAocL+u9IdonmF
DH6IcPogrCFPjkoRk3juirjPoz4IwN/hnuLycAcIKXPSi4iTgvsDmkaQs6GcEOZ0
8orpCJ0Kl7mC43NjzS9SVD8FdyT8RrZ0RuxvPmeV9wHe+eso7T371Oabo1CM5Uro
Q6rrAI9AUkYQDo1OXNfnoD8/pMnGXGnlSoewecMm9U6kOl12qsspq0zEK9j4GvHB
sJeOPUD3K0yMMpoSpBlxVbAERGbxWiHOuSRAVGsycNV24QkurY6nAI1X8WaR45he
KT6RK4DWI9WeQHPNq6M8uBY8J7IaYPix1njTJy52p4D7mzwvDr6cJ+ymI1towU7x
ynHwVwn/QP3weQ6EO/8IiwxCkQXlBT7yHZVPJ4f+xQLfM+v2RyxfGOAe6yYsfZTy
IfIxDEhyRm1ECYuTTh+UfZBhx2pQunqHdfvcXE3kq2FxV6/8qV8rSW4XU/bD+woO
kYzZ5hHa+TCz55HapPmuwi6+ZJQC8FVQ8o45TYsm3lb7Ls+9zYqhVvR5mcoJGvR2
fIC5wsBsloi9rse3No7K88hN8JpHKCHwlRBfJfmDbW2TMW6oVnlvRG1AOPTErs10
7vPZjpuD04HLBvNLMfPH6YntvStkn+rBz9PhVTYNvZnHaoW97ua/bL5RP7+EnREj
WUbLlrV+kl2duhrw/wvK433xzt6SxOz4iyQnNHbtE4qDXAggCkmRbdBIvEMIDssK
KHgMulMDCt8+nBonEJ5ImesC8egHRR7ZhS5Dy/2BIkBhSnmyvyuzy5ujGq0Ffoos
oRsOwRoHkKtWSiYPmrVyadua/LgmnBPKuXl2XGrBO4WZHnSXRir1jLlO786sxDDM
Zw0h/8DIYVUd+k3ERonoxOQUx7h2b3Sm8RuemUkEczP39u/e4p8kTWTSSdsmVt8S
I6nEz0Z4DbJpiFy7QCos2D3tF3iYeiXD7d4aM/vF+52ETD2pZw8vZXCwv4tCamx6
g+tFz57GHVSfk4lT7QZGAlCrn9NcC6xoFtVuIyGEYGLkMo1Z1QgkhfrJs+d5iOZY
QV1F0EwrAtJX2k6/MHkoJGBqfQoDOWp425yNgVTEw4XvuVube9+LIigGus41juj8
CBx3B5FnUP2DBM8pBzMHqzuQUfnmpMYA6ETe7Wb7idbvxo3FeKyu0PeYvR+7J/Wf
PIeE8cdlL15BspolHFQtPw8+2BKiPlkKCOAnUohutdK8ms3AoODHko0peBH7uQFN
ozs2+Dzzo6w6yG/T00rTX9tnD0esigZCpVmNn0b4IsDXOgyHqpjpN03tSgXkDBEr
oV0nFYGO5iH1zH+YjKlQnnXNvwjmTWvzmr3KeiP864gzabPWGHmydj5bOnqe5CDz
KFvIjy4DMeel0ccNimZCVQUSA7m4CN+X0LPwXxbh8jt2YWCIYWN+/1N8MaUfPDbe
ye79aIKEoql5Z9009RbXNRcmuxaaJSXudBJYc0sfGqFaEjIn3QHO9DWTH+rBAy78
sbMSs/MCu9NRwpEtiKpPgVVE58LL+ePrxQsUP+umFxB/oNGlUMdaCbhnMObJOLsD
rCVFLrr0wsaZCj8M5GhUWOERlc00sV0tsw6pQe5zlMFGkWeJEoP5KTHwSaIcjSVc
8h6EP8RkcsYKw2q+X7hmK16lbEf6U1MUDCOSjvuJMXUo9r76oKRTBfHpWp8IOlx4
M+5kILtVOS1iTezz/dNR1TUpCyUl1hRhbQHpM6xXJFoMCev3lpplvU6kDuEqkvS1
sjjy3+D+7aXmh5MXhd5saNYOQC22soZWAhYKynfMkonvmMeCVSNrxOOJsYuqN1R1
vzgA6QnxeZC6O1hEssI9Bq8XNQxSKE2JgJBj77nqzziYUI3GgqX9sL8eiojyDXSv
pTcJQer9g+pFTEc+eUI6VS6R8KSqdeughXQZm2XEj/dwse1j+lR3SjxTn5ipvw+Z
sEMuAekC3I0+9Mjqge2ZS+v/4BbFwkB8UGxAr+qpl0xZsqmM+NdGJH58qUSOP1oJ
mKR5uOWhO6CM6CNrY5VQh+2/sHtEoyOC19+1ao6qbRhDnIZQFvL8waL+JcNcefcD
njsxsdYkdfhEcJiy7Xu5SSHgGx3s12b7fAbZlbQ7v0VuFtKxCQA2CzYt+DQs054Q
5mAsjJ2EM3+F41PwGD2WIvEZuBNeO+nYNJvJN6NDbbh3hXXc1WPdRK7HE2pwat7o
NiYwdKnI2YLPsdfvfsgALNAQMvIQyyTzMpSq6tJNjAA8pzSV8kTk3mED/0l6NIgE
BmjrmNwPCn8PloBqW3MPTAU2YIi6XRFpfB/xzopbmBbX0oNbZZADRaBdfElg3DGA
OiysT1pSAu4D2LDqX/r8JxQ5PhMxYtdyBmTVw1bL2r1raTjiBmt6mN6QVOam1/Ej
S4OOquW3hewdgchYzqpBsGue65gusM6jNWgFD3oZ6L/xE1ZAdk0rwJ7/nMJx/oZz
SMjVpLsgoOQeUNKFDxS9hkD7OnWFC9naX2sJploiNjWuebeMrus9LNFmnfKwusNP
S6XAhT4DPmvG8gKbt8y3g3AfO4kLsZ2oSKWS+kBr21Dt30lqGGz7veRzqF1axjg8
pxvE9hO2O1COUj3xJLlTkzaj9p6FneWAOXU4zrOUDxhFiD4f6uN19+bI2hilh0tE
6lbYKufl6WF5dC8Sy255FAOh4lUC683h9O1JBCqvDnFMq97qrdxZ2ZHs6u72zMVx
YEjyUvDrgIGmXapNCSRfO8Wq6VhydKWNIVM2m2Xligwt6p2Aro5cgb3JcVjLjjyL
TUvUgQOr6Ho44Dc1M+mlRfuy6Irq8+ifV/6VSvpr/m97+oTwxfOxEjgBHwTtZ8/r
T0PVywV4kkmQ8GsCFCNdnnP6wX4uh7SoRbvnQyetZm9eVdVnY4ya7C/kEQm2XwjQ
4OuntAxUtEKV7fn2uAwluFDVSXZ7eUJ+MzXpADpkGzH6Y/qTqvpoQoLx4hJFPykt
pb1udOlAE5pFopndXe96kTvfSy3Cgs6znV/iIpiBkR95LojuwUgwx/ajahvogxs+
WthV0znWZSreju6Sdo+yasx4/qA//Lw3biuYfeOfKJDYm4cGmvzQYFQvhZ8BzOuG
9EHhsEnsh0zBnX5vpjZ5f7Ye45jGIOq/fvIud6DnSMaQcPOV8FhcDtdpTZen5ciG
+l6yiJaEypQ6d45wm7YReiFNwolQzoeJ1bDGk/VNWQzopWfkhA2gaEdmtgUBkmRz
+LBIOxElPrC01/5HyTi/5uzfwkzuRJm3iqavP3C+CTNPWiwscGGR7fLBGONxTz95
cupJahE9EtjetNtiTXLPytPBbBkSQBvA+I3E1mLpUfquWCbFFYidgFQJW2G+11xp
IW/riMGsgG1u49Y934MPKwsVH2CVTlw+6/9J9Bypp7AG61OJLtBe+DIf+c/4DURg
Y2aO7EFCiFmvW28UM0yn76SdHL7FHzVomq01oYCOmaZ7iq2jduQ+rWgP0M/RwK3i
fj0GwpDuxOLASlImphvezBiy8v1BopDLilg1quw1zOAk0jRGP1i9nzgxl5gM27xi
COTMQWi1i1eaCTxep5YKB7/cBOtXNTqa+QtsX5zBWPuYKo3GUnQcprFd1srbKB73
GvGhMrQIuv6iFecSq1eK69Rn6vmTFpnAyZ9+89hCoy2xjrE28YrREcb0pIaZTQIR
7ll1s4IkZIjvTVqy9Yy3kTLxpQKSRSzjdgM7/pz6orx1LIZrf06+l6i2U1K890dB
mR5y5pGRG+2DmZ12vpkZd7bL1RC2MHn5bay1q16skgKUw+M6E6HkxxFZVvrT1QRW
foUQm5Z7HRTpFWrVlhBH0MrlsuqlKuzci4ZNQqA07uolZ4NPRmHwBVbici0icqtq
t2MdFFMkrvt9FIfvvlhdDaEULgvojuM5PkANAZxReojONPPfxYVwD0cNjAAP6HzZ
a4+W9bS0syToiN5tDEVtHyStQWNg6dG7ri2UBY2scrTzIJKMghqsLFhEFM980KU9
PYLGieT81S8fNpKvtssw3zp/KjRp5MyGUBorXFyj5KzLOtkxHjyAl/d2FO7fqfjF
I+ofzg0Ikk7hSZvwS7hzHzxCfoBFqfUU5pWB7D5g8wV7VPh2MO8gegIwTiUyO9dX
ocdjtvZvY8CKNCVVkJlFkH9wnnm85388pkEigE0sHivjw4I7O6m33gKzh+XKMO0c
eiSBFyQwC416J/8aKyJQF4ITLiekX4+Q6GYCRsd3yWpt+bXlZhihFMUinq07LlVx
fpMbhAgD5sTf4oNkY5qSdaKSfNA2NimqnccQ+pYBy6zlIatkAaHrbAzAcnPgbFem
RFzgn7spXFBzBi7DqV+xezXVcr3CiN0KBh9rEVXn9EBMVBLB1uU0ZaYky3eKPK4V
kuhnx1fXF83uuTyfMM4uJZcz+ppkEaurGtKpJ8hgfyEs/DorUeWIAs/8123bjRbJ
MS/ACFX29mB/v32PRA/kGQhb8ULDGWdHmDEaFgBoevTg+RDuKbV9X7V6Jt2F3T7I
6BLnMV6DRwIVbLW0TSv/g2n2bejJQCsV2QsZyIyFEwBS0t0728vbm6NUgDKdt57r
4/riAxAuaBi7IJwtdDRKFU9gpNjpNN7wIM24Tr+9dp8mdmWae/B4ucsnK39iYhun
Z4mUlFtlSHfsy3WLPzFUc56QuxmeKKfYcxyQhTqM0ZMW6APDyBuLTC8wDFNqNUDi
Kf993AEe+jLAjAJQyrkIOgqF2c8r6x9adNOLxi78fX/UYGTbYTaETJR3W4IweoHA
2oA4v91haVTqOojWrIgR1kmkY73vgGYOmX1q1BiCAaDRJBGoiFh8TGcpqoZe/jjf
jV/eQ2OGdWg03UG6283j7tAyS5VTiAPQPRAqNwPWUvaea0sOlmEE2T+wuzn3N/do
eFu7sjEz/6NyDLFw1O/oqlMrdb70nT7YNukEBFYW2uOGOQThrGBpjC9eHY5H2Wr5
XHPWCpZFae+Sb70HknvK+ufYY8lSdVR5BIGkiKXpCm0Q0Z+HooF76RCSWH5bfgA7
cmQg7MbO7fysPTOSVDJ+pJw4ToEp6zDWjo9CSVcW7d/sixtthAztRKlzh2U2UkWe
B5I+wDP+Xh2ogHgJuZXaXxf/8nFmpG7PfsXuxcDsdilAq5frUG21w0u7+0hZjimu
vbWiuhT9dI0eGWbVOXjKgldgcYWUyuNdALD2HL64nm+Xkip969lVEzkjT2AHpkxp
1RFaHb+mhZihpF+3Suqw03yXNMnJtk9x1mtAJOTqhqAq49EYBESm3isX4yky6zWn
XW9GYd/h6vlSYaKOSJUAgeeu94V4mxugPHMEH5grOVOkYwMbNlXQHgrwe4gnGS4G
gbzcCB7LvdqR/baeHmmUPoI7OZ7pWyjH7AUCjBh8r1SySHUNrR1WTBHdknwYKjwA
P57X6lykktH2rHhtmUH+q71LWj+pEBTjDWP4yKqfZOiKMzkscPCiwVV5DRh4q7IF
dn+t7fz8QOCh4kiiXC/c9Gy8xZ4cHjoUrpBrugDaYmL6z4J2VcOGjQEhvbQJ7Rdm
elXsDY20MTBMRgFXIo52wr9jHhFSOxAQ9jD3vwD5CWqQdSLkpECacfcQ81QL1MYV
r2LLf0qDx3Vco6B/IMQo7AtJw3qaYjmQld7AJOUCahlTfvvOdRmz8CyaGfDHZ6NX
9w1plCPqDaO/WY2cyf+oKtB9BwytL5OcCpVW7TvOh2ZFU2XQkIJS+HUSlZd/jzOv
5o4JgXWP/26Q4mEHso5AZZ6kApw9IKkXK5GopJU3C1r767XeB6ttVnbvg1A5qVrn
zpFLZt2LA3JjZu8xJCgmq4nTlbOBK9e/Rdbxb9eQcWGoaa5jD6wZs9Nf0Bvle0Qv
Gs0L5P0DGReVtzVJZdeJEphtDYtLGbSZC1NqnM9HrYcXFthbhH0muomw+kj4jXyL
Dity+A3xcTmnOM5AE4QldBMcspi5j5ss2R/hZ+4PN0h5LcI7Xk6wR5peIR5IA8X/
4f42DHSmyegRmwtlht0RHH2jOJ1FpbHzghxU1tW+HU3/78LQQsCM9nWPteoA439y
QvI016GbttdXImhP94+7rZsSC61Inx8FsrW6pQ5wGS4dXYvy1zGitywn2B8UAddx
8UvgtHVUdRrSCABA8DIN4VUUux1rQs6RO9WeMG0/6ABaTMpmp2+9onpm8EKOt0Hi
uz781xQMYcmqakFMVZwX/WxsU1XDCWa/8t7mMOAEi7zZXUmF/EfZ4h7/w/PYBfxS
Em6Ec+Ij0nxJ4QBa8C60p79B/ROotiwQcxkVi4MyGXhPPGsTxA8iLBp2w6N9vj7n
+sbWMkmYUg+MDfjKMgwXoaC1YWiuVdWYeJf7i6MKj5Irw130FLrX8PIpXJJglFRB
euGsVtAWkDwuskHqluNsmF7XF6xSqXh1/iu4kmORMN5gzmhdQFFkmFFQHFnYu6QX
Oj2a2E6tM79fCYz+nh/qatoLVFMsbMaEhNyNG3qoi8vMBlZI7gMjhFjQ4kS/Xi4M
dTqSQ4Q7D1bAUswIwoBf1Jp39vYZg6B9XepmajWFIK+FwxE4eiJs3ackiK9iKYoB
UImpJX82yC6BY1TAwzckKBCIroFVZMzz0resKR+1wruO6f4ssz32D+8vJSVNtqsR
Fg7NC9b4BcwxggpwkeM7mg21XYdsEjM3QW+N7cBrbUP8mMnqB6VDFCRzz/ACzUD2
01NUlTS2F5mHuUPfD7f7XoFWH3z4LikpjLtTqnLoNgnVjD/52jefY7Bstg1vVCj3
9a4tGpn11FPtefHUpG0xyajrQBGxo7/ahBmgTEb3fjsT5h5edl6GM/fzC1dEY/oR
h8I3Oi2A5YbWJnP2qrA/rHTOq7lXiI4GXmj/4N+AZ3R2ZfLHXvXE9Fb8BT3FgJER
HhBUDMcBtPg9yu7c4bLh4l64rexePSQprPuURrnBsgat8YESRRnSynHV8Kj+Xvdo
Q4rof6BPerHlpHDcJ1tMlq8wZggt6balqXRFndrrJBlnML7FkuGlqZ22XIBJv7wP
FjcOhI4UOpwa4ozvxr4K8/iFsGolwIWaxySaVs1llS5YnQke+zjzyiGGv7DiUvfA
J8WreD/dJ995Zb/trQzGcB0+rsu2vQzNVNyGe2yx2mBse+jtpVlkUC/Gx0VnWduk
KHlye/PkyuFLQbUxrFiaAn78wIXlTXI4kalDnWu/wDm+3wlBdUNl8f1n4gRBZZXp
2Dkp9I3lDSEusZtjPZZ4x04Zus5twXP7kLPp3kyuIpcbp/7jAzbZPGM2zMDsyzQR
UQdh+l6jr2/z+gK9Fhmc20zRQUnPnZDIyBMqOVFyTFUor56d5UGDcXYe3EVCa8M2
Yd/WtL4gkpDBdHdquuyZg+D1FpigzE71TWFimTSeE8ellmeJb9JWZeGcP9NvqKDm
tO2dKxQYK5dsPSVFjW5cjQ9xdS1YQeT2hK7A5xoYgFmHaK8uduYKOoHvAc9pSKy7
QdUVl8fOKnKoSqX6K8RQLsQ2p/L4JS/RuK0iq162Hbp+ZMSeVDogJR5wmvpiWr54
xk8xmdjk/L6YzzAehhdc3KEj4sicUeivMNSzctTWzG8vPGpdb/W5x78aalUQFVoa
aMKLpoDWD9gAuMYR0bbOFhjkL4OieKSosuOkfm8P/B7HTaYzYwZrl81GBkc6ZjCr
Jc3ojyR0om8CRBaNq0u4viHu7FVJAtcFbk+VjgBQ+c1UVNo4/4af6Irqb0iLiHQu
QV8YODKx5YUEbcRKlvvmXn+NUeWegXGkDyo1KjJU4oGPwxJer5Rl2zst+yPzieZT
yOOiO6n9IEgSeJRHZ3EazHl8JX09A537l7xnccb1GpTE26hVpDnM4vP4R0JNT2g1
XJOKQ2FNqUkgRpxvE3aJTGImO2Eee4UCdiN/8QWL/2MyLCiQUFWl4TYarASivjSp
1MPnK2/Dpb/M4qRG1a5SqLc6NKwrZIOsmoYFMKb4W1gUy3xezdZhVv7/BDTyXrpj
7LdJLkM1UkcqAi6ybxZeVgxiR8HNWqrBtcPM0uncBOQ+MsxyyxL6NWb32TCoLsPt
IhZHrVwJ2ih4VmCotOmqBsLaU38Kma1fz8EG0MUfZAT0P5GbCd9JYgXuT3e8PYTT
OvGxVTM9EbmeCBbQtq+HQosJ3KsmCw5IITE+YLFZTTYW8M5JLqAaFI7gAkuozpVo
XtYeCzLE+aeQxDnT02jGB0zzhoADsiZTauClZkGe9bX7ERLi4sp9nj+tp6h9bVy0
ONB2mRAf8YdzdEEHihbe3WH0RpcyHaElgcKOd904FgFjIcumx3/9PGRdWghpJK3+
EdmqT/iGvxbUcir981XaQxkAavA4L5XywBNQEj7fPxc2FUtDteMf1U9C/Hn06/PB
ei2cMt8wqjfDmm7bg7T6+x2DGzLnYBFp8KajFnqcerXLaOtnncrVJjfy/e+59jsg
akm0xLi188d8dhh+XsD/MKW2Hw25jFF1xkw2tsqOx5thTaTrXkuz5dBeHjXj4fwj
TobkEZu8JgwK9+Et1Azt9LlOigVaIINoRVg+jNofaQO35vfGk5iBKiYNPz/p00fW
/S/mBugibsZKL4awP/XQnoCN1qdzci3ROMi4Q9tDCLs41yWerHhu9+subbD/cUub
YYj7Xf4airIqOM0h7gSp7TjbKIVJfKwRja/v9zQaydLR05HQuGWWMPDk/TBruRAe
u/3LfR5n5LNHLTBdGkdlZcNuBHDvKJRc3mY4F3/KEjLtMiEz4J1BY8o6lqaMzFGV
xeKk2N23ILQGf3eSqOkMsLBb5keebRX2CQjSS/7ZFdZfh+NyKb6ZQAZ5fDdR8tsy
D5jjjC1seEXUhZSAnb+KBUOa18FDeKG6jfNq25u9pZ/K6KqEdaAYGQA57xrsM2sS
ETxYnCw85nmE3gAWy+bayurRXfLYlmpRFcJkvU9LKu9o3I1SxRFjMdZ2Z/4sbzSt
+AwUn7j72qTq+72TYqcu5pKkdY7dLuEGyl64cjE7MTtxuMOFl8rFlUktv2Pqsvoc
ih86Yyec7cW3Fy+LNED0xXPybQ9xOe5wQ17IGmajUhbWO3DZzyZ50U4dYK2JJrzd
mgyJs3fPa/7Mk4SlQUlJNUBRCPNhRcqj3Uqt/snJGGVyN6TaIi+3r+sb3xgaDTRz
NRfnkq958DBoWLKL95pFL+raQU85OcHnMaMH4qMQFKrtSZVGMao55gLMW79AE7Ut
JCtYSWuVmxVMa6jskuP3sNvG0x4JXl2Gh1eJ6/XuOUKQUtGNCUb0+e2M/ysmEvg4
CCoIrU1HtDoIopBuM+rxtZAwvIFGOc/DlVX0BijnPVBfwKvQ4YAc2d8psL3omqgi
eL8u/+IXmJqR60cfMdG565GntL7XtCm79cjr44Jtij0UvIp35ULmOrPjxhQfjJ9L
kLVLl+C3HtffnIuF4O2z+hJtEYCFSqhP3h4tNOsKvOak2oBKaYaQ6c0RpY5UBG2o
XvcIfAlrzasDbOismGqSULoGydfB/Ylcj514B4WGsk7JsfNWoF0gZ7Og/w9jUVXR
xPzqlpx7a+zQgYfQ9tvZHFa2bgRY6mKxwXtsZ8rJUWymWNuQ2fSY8UDDKu7Ewj/d
XHKpABWwTszWcmvqicQi556JhOyMboSffAtLEch3SoVyLpYMAsb6cDIa8HsDmTCP
roxmyxZTtYJKmTBwKcSnUq20nrZ+byj9tOHD/QPNvgWH8R1dnTG6uVlxDsVnzpoJ
lCCQC2FFVllm5hd368qwj3voApMPUEj9Di9l4wcz2EPxcceS8C/gpwjeHBPMUdoU
sXo8YJ2TH/l16F7Uin2UA1/6UwQ9IeoM8m8qZ3QsB+Wiv0COKPz2f1d3s/HI4ZXT
T32TX9zXDwLLAGkQDDmgydxNhLB53O9ROxCqrXfrcNm1Z3zj8zUEojLM4cGr41qn
R4e1PBDCl2gsurMiU39T/BzxJRseHrfXWWuKs7crxDFOJSlkocr0AyJoJYtY2FlF
lKx9b7rzPKUSBqaTw2lKcdedNGFMOFxQj7TGxfGTrUYwchgivwRPrm1+pd4ywF0g
LFKHMCdWa/bQpgvxI2a1uxZVelSGHg0h1+M/txy+3Jj1CmSpZccVHWqkPMjc2f03
YTT2+YazRdR9h17W72y/sF9b7I2OLvDckdYfhxfTB9iwijj0OsMWvf97IeKPlRLK
fTBtIsIxoTNkrPELojCSO63YIILVkRUabHQN5aAFxQvNo1EOnxJOflv367bdwyJZ
qtTKI3C8+9TrbwXl434T/TUjnYSgesr5/x5tcsIDS8ApGKJfGGHpX7eUDNtIAaEQ
0DWnqiVM1/EYsPfVJEyrdf6gfydL+SzsdMdyUyucgF8YziGDaj8F/HE+bCavkCVK
y/uVKAylmJQCGY1wgxICkAYvWeDlXAZYYzg4oea6ZbXJqx8gEVzI+bbJO5RiMo3A
YNs5UsdMD370kZRez4dIoX89pDqHwunUrM4IOOJIq2CC2R6L/Z/LBr4EiaVgW/4l
VoenTqypTnMjZI6KhZk8CUtJ2/BM4ToIqe3P37JsMgOby5NAMOKsplJNZPMb5zYy
Hbpl7KdXh3VJLJitK+08cgZuv/uNcqh1kcmC7FkYsgn26ctbUP2jPUq6Xr9VwqJn
HQF8SwRDYLmIUHbIRg3YbYBnVflBLHcwhvHYUOBlcIQd/9lR2LsWUC4OIr+HMka/
D/hrmjIlVcN5GydNOKTpgxhmqc3FBHGS81bN40xISQzByaJefQRgrY+3C11/8cqw
onvPkx/9LuCHQv54NMIzNi7fa7djbfn8zWUqLzWxQl97rhm6r7C4pstpz8zeQtIf
tirdCrlaWtdXmoSsJvo/lMyD6UMwx05Aju7IgZaryai72ZoKuUBkyTWens3BUd5G
hgI0+101EvYh9QgJIMCR1GDH77S1f9EyM8pFBrHn4XCdCI9npANpTiUkFzYZE5M3
mV/6d6wRYDCmu6sBjjeIvWpbrSNKhBzxZuiUtsQlOxxZXGj1fu5PdLT2nkDl8IJ7
7h4vdlBffSoyVe1vYbC40U5bO5Ll447CxF5IUs0f4A8AWF9kQusi4EpknO3uZ9Ss
wDHKkxVkZXFKbbut9KAeF314j1OOEuNGNWY0FqaJZBZJ88L8YUKiarBfoRj8AvXS
JnAzK75u1Ddwc5O1xSgPn71NHrX79muLku6Khu3I8OkiVL3TBzEjubLiuPdSexp1
fshJWJ0X2koP619uoqqWkTupCtOZzjWUS6+kLSgErBgTyOG6MhMictyxtGjSmVVx
/DV6soO7rjZVQXQ1BJMeLFVpz1rHLFhk1E8qWo7P6n1HihOIOkbureGN0rwvazx1
PmgZDZlHoX5CIEB0DpBAqKS3T8/FLfDTiHnhAPeu7l51bMYb2wRu5Iklev5/qnU8
b98ZZv00czjQAcijiYpzmo7XaAKW4/Rc/BYamYaMSFk4WZnLx2bspkQJ/g1LFcDN
fZNQzKPRnKzroJ8FvoM73RhvA4HgFdv8X0Ec8hUn7GmKBbFjVoi1RyIc+iXePvVs
8edqg5kXUeh6dmGU7dWj33AhU4C16Xcbx8yCN3OYXIy2iZkeyQlKs0k/Uf4HVl88
Wi48TZzi3ayLfYZ/fySbS13OvVG1Rrh4rqJbKzx0JFIZVKs+uTWCGVSPnXmqSN9T
4AhKsqUanSgJnfuQI3VbUYfRnc32cAIBHWGJeBRUfoDKpARc5Sb3Wq8IFy23Alyj
AVqzo3bedw8UZjN+t3cdoSpKLoyfPOD97hf8//lWiWA0vZA7A4s6id5ddKCONiKj
CJouBgg2es4+gqggGcdkp13W7KlPo/ZufiUzQHcdTxaa5gk0bZR/WlW9vF7IK3iq
kHX9YCuU370YDB+MCxv7svmEHpoZkNnBcSokSIiwhOseAdCP+THCnVIr6vcEXbSD
+Qf78sVkLKQkZFpEUGzoyIYm1zQG1dEB4MdfDbjDCNzHxd1xFg1Qfpb7vQ/wSSdS
+YJ6/Gtpr9FQ+wAwcnsSNhPsXP1FhpWiXiZJJvXx7ZWtux/+rnCaRnjp+Dg7tjQ8
O2o2H/Qw6MyuLvoDSca2ulD+opWzfSG0NKhAiHaYPxhN18Wni5+xEWjv74ISnhRt
sSV3ukC3Eh6jbez9nQqbUwFQwrbPobCgr2HRxf4FgwQp9XZ+8LM+WGAclwcC6deV
loBhGO2lxXKG9qQLdDIn1x0HtptYkMK70jxTWilJMVWjRIlePtwT0CboTkH37ReN
QGcnlUXF92a6ja6uBgkaxPagRThPa5To7KC+c1bQbpnSev9OOjdmj0bIu8l/rUNf
sYO+OoTYpDkcLuU4XWsSqVaXVq/G1+IAE9na/+5Aqxux2yTEmfx2bkJtACcX6/on
OVp6csH964/9P+/sPKNuBEMLFwbtxfNjre7G4EM8Z4lFqvUf0BlvlpijdRhzh94Z
1BcjjT6xoKVXGAaWsNXWBQHN6GTorNPe4yuPcS966am34yy5vRq+1DwwjNiBh6i/
ChkEzIqLvcgF+PF+v8AO5mTb/b8aDZoWUfTPsi5JbyBIb8fS8VkUI8VpKmLvVkPx
s9iB/w5YqUkyq7LbLEHrJMcZcsmv/bcYPsxysLitE/zRXavf/KvJyFWcr4lLwVzl
gGc48v4tKvM6X6OwHYKdl3KwEjgxWFSijCoqvcE3958iAIXC1YcCNnJCQRiO8MJD
xisknys4M52h6BRm5+Bc1aqOg5kUKGIp76JtSrZCcDq1S3kvq4yMbpotD8pEpqVM
GZwbNZMbd8xEBwQv0fOIRMdIIsOyhaQbDat03jK7BhfcyYNsvJInTU+EdBGavoqg
69Vo7hllFCWdBVyDvuF3qazab2Ox78e85IZNQjBBHJESA8n+mVJjxVn1DNKuW3p+
pqm4nRMxJzE9qVcZ6d6kLe76JpEYcEmYcrJxZl2xGtCc8kqYOBWWOe5ILC57hk/c
2d74abezWXKOV4t9BUzZi/cPw6k2sWNSm1zLO2GuM4ebWzU6GFSUuntE7Dv+cSPp
cy0dq1HFsCfxHjanvTECruouReyaeg8xflHSkTS4gxDpPVFtJbgSdRXKYg9US3mZ
p2RTtryDhWcwRlG6NGNTgqvNWKTjGvyI5f4I+iwtROgw7xZgDg62CWFkbWIWBEu2
f8MnU415WjxdosdzlEph7I4UlyjZASvCNwuC+fkGuzwHErYoipiKWSOA5Oa9q1Yi
DAej9fMmFUMIAxkRClqiacXI90bIvGhk+IEjHw9NhlF2bDVZZqa9BMAIZ8lyD7jr
SCDrpa3thHnLSi4/9f5Mxo61mL8jQBAG5+SUqqEm0o87WFtaNrx9O6XHE/cjaNJK
yg+1CtJO457KGP6ceKwrt2Vz6Q43Wcspu3pz9mNo/VskaOMA3Z8ZlxcjsRhWseaF
IeAa2wppyEwDyutVzVQMU+c6AmhiOH3FG+QZJ+cjgPgHEGV8yV5h1sxpUOo3z5yQ
PGcVBFNMfbqcJ+7U3DVOKuaJVID2LxukZw5TaxCvNegda3WjiXh5QXsWMPleX5bx
51ODB1YQ2mVhLZBoItBdv8+tlKJtxCFY3dviBNkMWJSVGkHBU9RlYimSEijuc0Bw
TfpKKOXC8hK2vW2FaRA2elnl6vaLLi8Nhdy3QT9jMmXO8k4Le38s3Gf9a9QbY5SU
eLkUldSghdeOnEUVTJWTzJiNIcGZnB6Pde7Jg6LSBlgRWcisMDiEGuhaoHEDVE5M
sCg7WgkE4/+nPgOnsThfHerfcWRMaDumDXqMVoJlrArI+3rUFT1XNtNQqPDosVMF
6Dv8te5jqAu/5Z4ZWNIk9n03R7OeC6rwkLHJmXbt/owDIyV3ml/826yUcGI/RmDO
fTrCsVHnEylKulfmP+BxCKV7m9vcCyQpw4wRGvDD8pg/e9Q40stGp5nyELXTnivi
+Vgdrg+Th93I1I7tHN+yKLZOVnf+GMINAG4mqVWZYfAGLVS1pOOuKIkDJ2F6whSH
BF9aYHkQp62++qtszmZOVLN+fx8GBGfK56dgMi/AhDmfb5WEgovOoc4pbyCvTM83
GQtB+ZRULijRw1g8zsdvzNXiHdqlpZrS1T62yZKAv/yYWxAw5scmzfrKuVc/dXCZ
egdOb8UHPN+WxaReHcvJxYvcS+/RHNlCWHA2CUTZt5UZp6BllPQnhHaCa1kIiHye
faGdOh50oChwwZve5kvLzT9qMW+KmnnsG4I8Jll5p8Sq17NOUajqpQSG53Ijh44a
o5jQYWRJ43yxf4vfgxeVPghnkvO2g4VXzB3m395lAGnEWHzD441Y013Luh0vqOnx
o6HjwEs91g8VUOKQVgJj6wSQM+4dhCivEIsBTvvEUmqsbCFGLNdDs1FUnM/tUglv
UyupTfmyspXVaKcnlYZ0r+xYfAHA9dMu7vgTT/evifD1hpP4Bnp8tkX5o2KlNm3i
F6YgmzcihfTkHZQuiFh1LhFWuo7RzJg/kvmgMA+qKJfYYvTua2RjqNAWZs4lOMp/
O+goD2mLjxnByymCW0KpP6j7dwlNAFRQi5YNqyVlquol3WINEtVg0kAyppF/fII+
LgXJ8k9j/8cB9lhNLKUlZvmn1Dxomc21JGQtan3pA9nAQKRvn0k2VU8CCaVBiMtF
DF16zCzuDFSvdvQVUqaIIlhSC01jYhKAA08iAVoF6DFXOToIKOG6jXznYXeblMeH
GS8/h9oyBsBAaUGu3H75an58Z57zuPdXYX6QGxoEihx84soJ5tD1kxFYPbBu4Emd
7uJ9rK9ZPOziPTAkJT7jS711S1kX7FilFNgg48QXeBCZndiRMfwqBCuQX8bUSLZ9
cMEmJmN8Jw3PiVXGmzy/3He4FiVvh7Wd9iudXwtpfRxezub0ZFhJwCgMCHLYoG+V
DwvPuKdDZH8am6e97grWPEY0PRFEZzjj6um6xEqs7wQTzXrzKvHckqvksE3oPGXO
dxejuT1AeuuVpBn7rGYtaV4WH3iuOn48yoWk30HIh0rD2qmAJ4C8B3KD972FxmCD
1e/fMBdNiFPfQoBNks3cpNM3oc0LCOI5hR+LaO6/BLvqCnXswHWco7JznjG3pVLs
aqkbMrxnuLpWpbC8z+JPEwL42bRTLnf6rVaT8TdIwB0xOUPIdKnkHQIv9wqPEmtv
N3rJ/l9Wpq4TW+1O7RG2RsSMWI0uo7XeT9K0pvN8U2mgcUXDpca0C/yhK5VRnv9/
GIfamhdVLE4u9Ufy19ZImHVqSBHEr3IPE1I3uLPqlgz1+93i5LsQi07l65Scj7gn
7M3xRsMc9KBxODnmKe5hzfGHpytN3JAo9v2LY04uhhA0mXQBCdrHi34WOtQJBYi2
BmFdo1zAmqa3+yQ+ApsK4ittBpuToc8Ql+5SCvjnKFdw3P1oOuUk0tKtMys+vCqO
qo8HApK6dn1d6dCrTni18Cas1aUMzuoAaGABnDQFNI/F/5OTMzGPR2u9qFt9SuC+
Iq6pTmNyNHjBrFuDL3LFrcntPFe4/Ybxno8OLLmU+3XBLPAo2Fi5rfnQb15LW/L8
/XvZ6LW63ilVk0c62wcyViR2rcZpCDxT3KCA6OPUJy6CuJs3iHSDCBHEEoDN3KOe
92KLxselZwfAA8cIfkLDDz6JwUiosOeQtvfsBcTbc/jyDfL48G4Anu8AkVYx8Xvc
BYzxkA5VrCL5R11L0PExWYkkyin+jYZhBg/Ug8GOWfsiborBxyXVgF3F7ZFgBDNU
ym3aNGLsAXBWc2KwT3UmSxYh3O4SUUha7mlYP0lUqYL3VrN6/GXMM2CCkPcHrua3
s0uEKcs5lzzlJF/ExqAH/MQVj4jt4UGcC1DCecZFMOkubULdkdDAfVv//wDV9HAL
LQqlk9jtUNC2nImGkonNuv8H3PCEBcEUCIvAt6qJ+BhQkLlOtcXvAt3Dz02PrN2u
dOYVwA8je8zEF7IUPaJggTJK75hLrkgv5DWOD5r8cPf+r+fv4viO98JADxgXjljX
fqXZ7soMdyJ2cxxb3Zph7e9eJQaZcZ7Gij+xsASV06YMxXAvEIFLXFOp52qwF7nY
jNBk2a41yFvXm937BzVNdJbx4pHibFVJAjaYagtm3JZxIaGbO4wzxbHYvAG8iHfC
mi3MpQxWB42VCopY3uHoNPOyUEutN3uW5vwvEeQmyi1l3sqE8OwcfrkZnCwqqH2y
V64n0265o+fOK8mUY1Ja2GLe/9DaE1TNoMVJeGi1SnZsKWK1QEby4BTAtMmz6HE/
5R9sswfZiiSN93UleZtIfdcAlwt7whNjqgfHjYcbxzFjEkU1tJ/usEWrruX9MhC2
nIJvVynpW0zBBzmn1xn5Z/8YEZIRVaBVm8zyGXiKooAOJkEWxV1MDSEaGPYqsAv9
R6Doo5v5wWrFFYOzNFXvqR/mACd5ZFRzD/wDCwE0SFTGNAHNuZn7OLKCk6QZA5PG
HopthYnP15I5Wez46cDZKOmsND64iYVt9ch/n/OB+Y171/zALNYacGyFNnlQpVF3
EWLqUYu7usn0qwKILD7DXatoBO1PypvVF4ghApRt85H/6GNSz5Ku3XN+pWNz+fQ1
pj5KCpvTMImazcCaSI4IDpbPK1sqYDynUa8OHT1cTLw9w1wzAF26frtURZFiBsFz
2N1AfCFRcbhQ1s45/ssgZD8Rb3KK8s+awTejgC76QNimRz+Jwwl09Aq2iap/+HvS
SINBw/RT2DI814tiz1xGVwNUTsWvE1r7O3hYYyie74tgVpzChhme4biobGfWSAqR
wPtW9OhPQRGzkxmOHlYr1Uiv+j5qWy4AGkAdFg6z0pVOThbzIbWtkxpOn5pytwpF
NrPvsTcOcx29bVgT2XITLPNvA9b3aTbfv/45abmAzGM9GAWqOEioo0wOb1pTy09O
Tf3Ns0cndCEbw+28Qp883r1KnieFruVQRzRaO33tYj49n17x/cKGh1PtWDzX8k5S
2sWuNJMQ5dmQcp1TgnOj2xcCyGYPpO+wte79fl31CMkaRimN8dHLrfvFK9KatKVX
YnGgI+Xo5HAFcvjlFdbtvKzRkYRDovhP08zHSnpkxkdlnyuBjqeKuq5X81tTjNbr
GSdsZ4g21H1nkrK+t1PV2P1fvKB9Q4m8sKBUwc2bLN3lsfDmQ9Sdkw5LlHI1N6oq
6RJMzuquRAO9Tm08bcVckmvlUocSS/+/IwUOivZSTWQWoLkqPES47NTBFM/fk3iv
EHJDc9Q6c1fAXLOp0N8AK9+/dv/7wlyTWNd+LjnSm6mrgiTs6trR6OjgGSZmWfB0
UtbQZZ3nBrVb9/ebQFoR1IYVZlhhjqG0moOl2KscEq14RUrEAe+LUf2X/xmKPgdw
7Bddoe0Xe8J6TXAmEoFjtyRk8rwmaevitlDwrLIK03TK8xr1RZYmNf5LXrQyj3+I
jTcdcKe2NNSFVpn8gfeZSD1zCgqpKPHn1GkOScWH2lRSU3kx5S8mfCXOyHwSD+dg
+fUU4SsrNpToOYPxXU0hyubXbl/fEFfn3UZm2o0JwVv1bhYKoTiMpHLpLGyQpSpU
1IYn8VsFdFsnNCvUOnTxFm4qYACSwr6Z+FsD6JW09U9bSR6a5wK5g3D0xeFjX0Jl
FATSzgm4AcMCpwslCMv+y0FjVAJY5/fqAX5s60PTvddHRiwF8Upw1dOhw9nhtQWr
ROumebQSgG1jjAmb/bSX7lbDlcS5ndy3kQvMA8Fhj1wR+kihlz4tQsQs9hBS7TnG
DGIbDXYrPXXMCxhHoEGcm0z2wDgbEH0JQizZHarVbUh7FXFonDb2C2U6fzVnPRT+
m8aoPMgb7BvcptCVebDayY2p5EiBDNIW/2398c2myznAhY1n/OC22Ed3eK20dOY0
6RHLJv2Cckposvn6JZ44m2X49f+mfH+MaKsA4YSL+5RJkHR4mL8YSd8oYTsAbu8Y
YcrevN0zkI6Yo14Qfxvbt4baoI1H2SfGApWI/DmEBLZlad91oQGlFh9uJPADv+25
8X6UFUdf4gt4umxFu++L5teZiZ7QPMCrj/MmB6ydiQIxUB9rY1uSpMBE58M/xDi1
ykCuut7qeaFB9JYZ2Dyh/9ub07kslmoSMfpFlpp8eiPksEHnf2uaQOVXxBfya0iW
oCtkJKzus7D+/L4TDaZkkQyQvGSfEhTN2/inYtWpC6rtWJltH/YZr9QrUgmklY5C
m13cZbzeKDSPZs7ocKv7QHiPY7pS2guQwh3LpAboQK6Wnv1oVmN0qix5N9fPePu8
k2QcjtAdVfFat7Zmc7y1B9xDWTujEvA9+eR9HEdOQFAt4+Lay88tB5k7cMxz2eCS
D4WkQsLtjfm07HAdNvUZS5hCMvciVLkz+lCKAU1DhvrxlJniMqTB9kL6RgBxPjfS
nnm5wsgcEjBcNoBdGp3/8iofUlkwj9wcT0s0Ox8kiAelTFJdUqSb7OSgFgL5KSIW
YM4iVZsiZFBkZMWv1IHfCAShCcX9twsK9E2rduBoVkenMm+pJwhKEfUmWFIjjdST
XgnLaoxBtZt5Be2ZDcM2DgrU4eXEPc5E22aSCCnaM4RwOJ/McLUhMZ2I+BQc3aQg
FccmiRwRgstEufCnd/9dQ8xFd4RY1O76rZ0/I6bmUJlKjvBal7nhHDHqPs6d6W6F
XB5SVhLIwC+tPzwLGmxNN1+14DWY3xcIPilAG9sAKFl+lkSlrJqwMXW0/WqFvE55
sgCTgk9DZX2qEW3X+6vHP21kowOl4oOwcfhXLCIAIZOb3jvU/AHbWUopqLPW2hgq
wY83kBVoTj5QwN18RBjrirGJ+vYeZqMCSObV2QbH2XIu1lmOfVkZLkBn6aZERhGb
O+yRWUEILKqSHlnM3Mlh2bLRAPCfPXL9bx2WdUB+W7q/652H4MUn8dyz8pmT9H/o
ywFkfuN0Lc5RUaJpLi52kyPGeTONnmr8BEbfN2D3NCvXL9wip/8a3+qhLsQNJHs5
Ifk0VDIvmlR/QJYte80CffZdncFioll/5saYqjXg6A44Y7xPakF6e1agjkvMHoi7
MNtlrwI+EnLLVpkjbK79CwKFyN2lI1UDW1NxDnoOOEGLCv8fyEN3P8JurOxtp9Kx
EFR+TaZ8AGMP/+vBCClfcMemYgLG9yiemKXl7pa2MjDecC5tgQqIksUOGCBsjJz1
BFLiUlFB9WFtitoRn9MpYFEF1FuJQCDuUbRgLXWVEMps0LL5J5CPuv3muWfFcTnQ
tK0LG3UOHlDs+DbwTf/60zbHz04mqMxH48u4Cj8YKGJE1OEuebO5upcHcSYNYRN2
SjAUPsnOLpIiW4tbyh+OMuI9LCImUucDIgmXhd7LYYTt5LU4dKeN2DHwyYe1+fbj
oA+b31GUktVjHpXohRfA0PIAxCW4I/uQdyFDmRg6IgA40W3RKVB27S/F5qOnUmnb
BRcyMZgfY+lt2clLNl4s+7uGNn5Bk1EaN7uNLrKnCau71lDLRqi4H6SMfzNbCAOn
YmPCE9p1zLY1GcTmcKkPClMOL9V3sfHzrKJ1mH1gBuo3sMXDjQ/PQaASt7Up+HUh
8MR//XBvdOUb5KpiMXsHxUWjTSOaHptFAgHfUhbmyTEy/2bpwOokHYOWcdITR/Mu
8gzMMyS04MsJQz5qanIbAEgbfJRC4ZfCq/L8v6rIUdV/d2lkY0Ywpe8OVip/hlHd
8oQz+I0XURyGxI+epnLGF+KL4bJvp0jIkpZCFjogJYBW6onmcaT9sLueoR55XK1Z
wGTTzIZzMm550WMljqGY21pmkL2/WSKirC97G0Ajaz6DCcQwIQDcMiwWG6S5bmX2
wLwlXp6/pQIDdAucgFudjdHETYDXcCm+6FXuXf2krXJyi7hd5PLgsj2yj2RKrT8H
dOcYgQhyixX+aiNFZ0JhlB8FqcqbXN3BUQoK+FqxmP0Dqo4uZ8z2/FJTbk3YUfUF
25UDZWIoi+hZLB2oPdD8+n0heJAuMd7vWSIyqzQzeK6ijCTyELrfNQwevMY7guB6
9J9Uh16sTnf+x8hw2VBP4FeozfoNskZpA5iUD/eHXi8zdlloSPA9PFksz7NQmdYf
j1FGDd2Wcmq/d1T1YDXibtZ8nAwHe8F9ipVZ+3rE8VT5+6aMLp8nGod3N9go8pUH
wzTKy9Agt1lfKdo6F8etVphhVMcl/7mUUx+yuXRmJ3DGnOYSwqWdlLx11VFNdx0U
z873hi7AhjITNqGdL/rovQxbYtxg/uLJn1DnZGU9/44WW1d4CuyVdhRPJP1kFh1N
o9UD6jpFDGL2KC/8+Ey2Gto46NNkcYBIMBwf+SlbcIVu6sJ9tftpR6osirH3W5lG
nocxOpKRWv8crogbKpjDzUh08/lmfvs9vbLPFF63Yg2tpnKqbpCbEJNVMOfnX5A2
om+BF8GhaXQjs7NQgt/TH1ZbLedW+H4nca8+UDQjJHI201eGypKlrAIJDRIdOgz+
q4gbO/s9h4F1XxxHERkikoZbwDQTX5loKwEzBgsyBIFGbkX6kOGfxcVNGglOu8oZ
Mald/Po95jLi0nDPtoNNViraW5FChw8Y1QAwl144ks02lpiDQnwHVcUmipd2UQMC
wrfegte/1ee+RtihexNGFQrMD3J57ohY+ZJ/AwKErftSQJqjsr79yWz2tOGX3DwH
IRUA/vxzR9soGbcg7E829+3HdqGDG/x8Nl8UZlUZjsXevxAiXPX3p9RybgvDk1cn
g4d0in3AATgjKL2T98Inf0K0zG4bKG2mHLS0n2s2/O3MBHrLN8Ny1dCThIErtnAQ
Seu8sLwO1hvNxXzrXoG5NYErKN3Pi6F7d0uZjTaKcGcAXFUAEn4/kIZAyd6HACY2
F0de3FBk9qHSlPgtITcbgvIGvCsyk/AN05FhHNVtqVqRXWxWxUpwIj1GhSTuQkXu
vmd8+nZTzYvHhM2swnIyj2QqL1OPiHBPzhRbq1qb0XQN76t6S7S+cQ1w7XUkCZgF
K6sOCEhPM99dRFJS09M2vZWkLqNbkPYOfO5D8NIqwpUkqJ8C0BiiDvsrRCPVi9dy
pkRi8bHEL0iIm48fLR/CRm88q05ooZOP6aFKAAsWoqO/6BXzr8j5ZQnEwCpKDdN/
MNwRQrl94/7iu5+pjbe4xySxZ/Uq+UJssqoHpjn2Nj0XlVHoNxpTLSepp4o4rnDV
nxzN5MEdT/qvkK/CQP0d5YoUFY0CcjLG08COVcTcf3uLyVKe9MB8NWLf7XPE52Ex
2Qnxb1T5OvdJJfNe+XG+yxko5DBHOfs35RVuJMCmfZo33WEa1je2Qm+9+6vk9DTx
Z2ZpAlw7C5QlW6/71Jthq6NuRELGxikovzF7fBssn0BgEGrAWhnuGZgSd/qatAY7
evrWmnXIDZqCtQVP5LbVzki6HXZFG/DiLLLNnlMbbBB07V8EU/XxEBbeQ9mOYzWt
hFzmEpSdT2a/MkQuSDkdQjGZVlDb1LzL3BzLFV6yZZsDYIl0EG3iLjD1Rcme/bUr
V4oeuAeDlmYP0PIaqTk/ozbwkAoF0DQIa8eBBp8rn2qXF4gQIKHij+V8xCgorRoS
/pPL3+/iTnEvOr4IuKSJIIpJpOv/uhm/jiRt6ztWpkZhNLr6B43YJj8nWgdqNLWz
875ou0hiS//auvniAj5Oxb/zVRIsiNPGjLK207ZwDnmVFLhz8rcV8ETnGfwdKqQW
dxGfkQ17tkJCIsI0P7Ckk2iPpLIET4f9rJwjY2X+WHb+OxZWjUj6pxOIXECOr5d9
4xqTPzfVLFM0tuwXFWcDZcVCqlohDgp0KxkT4cFu5SAsXDVo5NJ6Xw4kz0FlHemw
R/HDJUQkj3b0dosO16Mwr6i5U4y0wbzwXlkp5/EgFaeL8xV1Po9cTZxkDFbkPwl/
VAhbnzi2FdwL/7EkTZVcUelFGn8pbJL8V89EZVraD/86sGnBEiKGHYRpLgOmvtAD
yT4cncsTQ1YrbxbdeVe3I6EBw50lmkZbBjCSsVS1YVQb+N1HhIagG2sSsHeyfoOv
MCmrR8uaooxc60zzU4ihr6rOjB+zxJRifT9EM2uLuZ2a6YhQpZEJk9xfms46+b10
3vB5knx7NoLhZA9hugDiql7Pxhg2a7GnYFzrHuc6iWivS1dcki6EEuiUA29Swr4N
WvopnkYg64JDkX4pqUfzWTYqoqUQixGGtMwYwQRReXPipkCZk3Q37GmWysHDk29G
LUtOSE7yCCR66unZuy7NwGSZTTgE4IaigMkU2Osb1hSBdm1p8BwtIYXfxjY3gsbb
9mw95+wTs24Q1EH2MPMEwKn2ItBllomGFPqj44xsf6hRWc2bd79FFMTurwoD+o4H
e7XQy9pcECcmIrpoR+shPXbNj+fX1qJYRtDgAhsfrntG59s2CF4qaxgeGkCTlPut
0MHgJ6v5xIZA8VlcqaiargymquhYFjZ8yViDW6pJxDtGMiBJzeHqS6fdN1J1Ga+w
W6CMqlUiEiiuF+x5SUikx3qkOqri4T+jBJ0wGW8sVLGgXzYq2vnpEN8mezMgaSS2
bXkyjvphZFjIrBPpZ2GYtRLyPFvexXvjML+dq1oafqrba7lH5P3Q/vSacSJ6Uqyh
khEtz1wm6/Sh6qYXo3Ybo7JTB6dh3dJUhrkUl7XgbwUfmcxcj0WK9ccxMpet6MkG
X72zI8ZxLV8akDnTLoNCie7HXl5jo6U4WUl5BxFjd3xEP6ra/exsSQwT/uL7cZgT
u996KB+Yyfzf6qi9xdzPNXNa7d8FW81zisOtxPwGrlXB+mBDQXh8deki/TAAxp7N
hevuJl2xLzGSlFdeSkqWuT4DL9aAsI1iAH9iYbNXA3nSIbhAl4ROyoiZZG5jliuw
LVgcd120X8Go3ZclEp2MBgMhaw7lzyFnsAjHaPM5jHl69ddVn4vOmMJJI9DPmqZh
ac1eryGyS6PrZRCw9er8igUuLHvr5rl+dF4OtsXZXps8x9CwSjcNdF/iJ7hPqY32
f6K2ReFBoGlAR3ECgTyFjS5HLV23Q6DLJPMV+yCpALeuDo64RjhGOrBz5YGXvYZs
KJFRC/VWgvFvkXibv8FuNSFLjZJVdPGrxwgYkEeCToDAI2Rssq/+QtcAyONhzfvo
fpVX16BSYavWCqMEltnPZ4wk8j6fc2QHsxR1ltNM9PDYWZuyTsbAR+/sGNAlkMm+
np7T2X+tSSb3VCKOQi0WKuXGvneVhGW5vRkl786zPAN8KK+3liMBNecZV2fEzE/O
UVWFvtWOPuYIXLCcrnPzbWog4zpouOHi2xr40s7/66Vp487qvuxQJThrmIw3I08h
r6WJ7Cf5tU+Ij4qyPPi8zEE2xqMtCEE210qwJo+eTPslUCiWiBYO9qrAJnGo2qd4
MopqWKp6+sLngV5U6voNFYHRnIY7ZRV4spcDSyQEE7AEW4WqEpR4G6wPnfraD6MD
EIjECTs9i40wkCnldWxgJeU2Ci39MTsyT4UXEP4InU3BOS2vxdUShenUt51bmcFA
d4donirPTWN6G9yTjS5MeshYHZ1b7bKwLOi8p6AsVytcTT8d9VpqXrHm9iPx8EHs
qSOvpZAmgU83x7zYvihAgmxyyQy6ety6RjctEAPf72PLactPGgEDKSJ9DUgH/DWk
dZ4vmlq6qmEvcoAax9Vwf3UXCogiRTlA4c+5xKNAn5jrgQ5UADI/yf1kc5SO0Msv
Gf8HJkdVwro6Q0og0CyxuzCebgUJ62i8GbEZm1kQVOowx9SNVKyZXc5G1xmMmQ86
zDiGSn3CtG6VaJBKeqrdY0UTQzW+Y9OuqY3mY7Sikf3Z5AGjwV95XaxU4kexY+0h
4qnAdjZJ8dXmOKXnijX+A7kcGTFwbfTPieDK1xMj5rcbWUJW+2ZKPjLTCPqhVpo5
X7Rt/9wxYBtXXYduRGrwF5XNU4TqcfLBKVIKuQ/1n/nzFU1nND3ezk4OvW0MwC3P
f5phcHbkby//DAQgCeK8fi+BhJULWMifGBA0IgLKlf7UdQgyVOS0nj5GTmfr6WPq
SEjbgLFbrNwLn29eazWvbvYqGb5ledpFx3VCwwtL4Du5ufjf1ubLLye+l+TEWpTO
/8QovEG2Ip9oBzUSVxm4HTv1LRsrznSVVMW4Ra3vdrgPEDhi36UtggCjq7KFPRyx
C/QKyqFKBCp3/dAKwDfin/sBDHdY0OHMgcGljbiBbxUL+Dvay6Z0knLhGm8UHtOR
Hazci+DXNHOlR6rBC0wfe+vWHXaiNdQqL4PZ2E9ztbYvnsVhoIbteWyBE3q7T1ZF
v2eSNHzapFBPqxya+2BD4SNokzTve+H1VPeXpikK0ESouT5FRbs+J6orUR6jAq8v
Lke3Sw/dXpBm9CVkyPIMCjigcJQ7LFa5YQo+C7DxXSvvw2CuQruzNsx/c5Ein1Zq
dby8n7EQ4S5pyYNqrkjd7X/bdqJvqvh4bRUJP6RvHHk7+JWZ3rVZMANdY9ymgX5D
ybidX3swzdYAM5I1gn+m2rBAWi+rYpEiikVxQceF9akt0O3Dy+Uje3zJopfgvvZ5
O5tGa2ypUfFaeX8zxQvaPygPdkCIj5BrzAGoAqxg+y6XFBhb2e/L3V2R0gAHif1T
5bB771CwyrEzVhLGte2Vu6Vxk8Bx3ikNKMTH3Z78+mf6vJM3n5t8hvUzZDFwX9wV
0nw5JgbdQqyl4ljPWnkwVgE5LnInVxZDZ5Uz4mYq5AXBds3pFO/X1oznx7iufwlx
ZB7ECSY5SqcPqQI+bX0UL6BmijBFwmbV24mROu+hfujRNUtXUfEJKMUXPcaxWxJk
KDMgU5Av24uqqmiVvCQC8RIZvTFyKUFdfXmtOzdJtdMkE2K+EHZUo2X6jQBL3B8X
QnsZI6rdMaUVMATi43n60JY7ZrhNG9xj0gF9Op0n7WpwYVfPlzJBiBXsOppUPCcf
wNJ8vG+9GJ8S/0Y6+N/O3xkb8mBqD4sNAegIOvo6UwKcgxl5mh1Ikl/gAc5ElSb+
3GPXaFIfCLbXS8kXqhqj43tsaDC242gvYSjmKgr7Ytm7UsUwq7+90U4MHTYAF40u
9mvp3PAiGJARccw8CMn4O4WXj+VI+nDsOREZikpbfiV42RqV0ylNtjDNTXDvndfG
wVbWagC8GPNMdnzggdHIxBUIcVf0NBRQEdGVyeK2LeLW3UPFanAh0UHXXVUmVr12
6DYkyH1SpNOW5vqukBNI+xtIT2bNUoXXezRyt3A0r9JcvRBYPcbq9E7KjlQoYeDh
DYscqwCcJ+/+510eDekmdmHhYE7YY88N9T3/LxgkvTMBrSuB0jgb85si5iVxxt/E
OVAIvAvv+ucuIYPOTV0GUkwvDmDgj1NaFuzaFyktdmp4CqaPf6VF+DHF0uVogHWC
DI4yqaPpyYRNlAKHlDVNTvK4pSOkcVnFCLt3LjzVKdSOhXCXuYXYEw+rO5ft+jl8
6Vw+/0+yiP2mbnQi69tGn+t2Ru0Tjmb1QBAjYWQ7EYPbyPEMIJYBL+RcIPjZdTlR
a7jhmILj047qky5GCkhYxF1SqDQS9oHcuWimqJpMClTplcrUFUrJcOr/hTQJbdEI
5Vj/irvfyMjHvMwKb7uv26mrZnIeW9XyREr88IxPkRNfSC7QDG+U8/jnECZ33FsN
1SYQHU8LMlOYEzh+7dRMAQwYYZ7HNa4DaSuhhLnmAki+N+Ts/iN5ZU3wsCcHi6Kk
OOgkOB5SGZ3J4wK/MVcSuZB38lggS0PoRAdcHLYyJ8yqWA2E8l/Sp33vykq26ukG
IXJHNABvlS7l3YfjhMirWVsky7OXsR8dL2DQSGnD8UASCijVeYaNHiCDuszpa0UH
k34yFp3v+vtIyHtdSAQexr3cnHY0T+NwzfiBNhwqQS4+vYPYQYQu0zglaLSRUi1m
UVq7mHKaXMkpRUq/U/IqACDsQ0GwkwD5XNAFOyxWFIhkoC4sUS6seZo0IbvRrM19
aa5Vse5wbQzdmAgl0N0pYyYUHjVDjlFaBsyAGx70r6qcaARtBLzcITS+HwsED8P/
swwsAqDfbBiJQmlqCU6SIuji5e1+cQMxmeS2p3HEFVHRKGK3Q5rLvh31fwmT93/7
wLucuWBd0op2QlN7MJ2m0qeiu4q37xl3m3El8sPC/5CWAqM1vjvvnX+eenJU/oa+
b3VR9Ue84SrcY9sIGJ8Uep1bXdQmsyCID0qzN4AEiYfx+ArDhJFBCTnxbxJ3xDBV
4C04E1CsUpWGA5lTtV7RBn0knSmvvoAKGnSoJuYnXwlA+md/Iwhq3ptpUJkPe4QA
ZyD3fdtJw5kon5t6wf1snbh0e4FWK2esfZ9RvCPZ+ebZeEffZlHHgq1zRBzIAFYa
7ZMAho2Gfl34bm4QHGcY9ueR7yeL43hwBDWiAWTrjPujn4PPahrpjfgHj00GbzV+
ESLoFQmSyFamNMtDTYpZkT6tYkAbMUiW7Yj0Mm+giRE1v+KpRACEOvoITnQP+p2g
hOVf/TbN9RtJCqvt1MaeAvByMEnfidVYfFV81wqHUHf9m16iCpk3WmAZTrOgDi3p
uMeAL9PDviur5SyKYvcH4ffSAwTPKpidv55t36A34TV0/B1wvbxxU9V166KrZUe2
EtYXLM1fZcZjNTbvL081T9PxsMIqpaQp3HlAschso/EP73haEAWZXdIZD5IsFGfV
VfWMzjEYXeYyiOPAt7DVI+vwE2o+DW2AJOqbEv5e5nMDakFWRpQrjVAoNuOb6mfk
jKf68rRsLEWRQK1+RCAohEKd2PwKrjmKa8CU5ed/qtEW+/MCuWndfHnEWwjsy3jD
GIvlSQfa9C637jj1iBQEJ6ez0IF5KknKRAyVvkSmfCGIFNbm09IkM6xCqYnBVzSc
RXYAxDG9zk/6umRsnY4krPLYZCivHJJqBP3DiRxryZKVef3TQPpYTRpx2OlOj7+a
5qmTJryeUrdHrrHVW5tFH367niDIfb5jVFvDB19Zvlg3k5PvwdrqL8s2Nmh92kvU
6t7LHyejik/OminECiBwCgaXjbyDDp/jQ0uZnbe9LD+wh8FlqZFCu6ag4Hzvq2Lv
jcYIUeyhzyyUJzdBqyUtYGGKuM0KIzS57PpykARcWJCq489ueQzb7lgsbJyqjNll
jp8RtcTBdE8jX/MaIFMN0/GGq3wQPcU2jLSKDkgLW0xb3DoO3CU+Q8LJYCPYd6AF
5Yd9IeWBh6YCYnmlKhoZz4bkaWFAyu5ff6KvG/6dHx8nGOnAGR5EcwUQnIyGmCWr
yFGA0IZTQR43i5RMexcqdrhixAtmxBN60HgxbcSrmWt3kzeGW+u+yhvIwsGaYAGw
5oVB/F1XYT3TE8xxahTidpgCle5a0Lu5DOMvchAsg6udEEtU9u6prgtHUiirhSov
xEpf3kd4E9aPNdoYg+hOap7asrB7pwhiVcVFMixA7Xv0H7wIDzWOSUMmzaqdWQfe
Qb+Gvaln8slIxWpYu9jGEXEcF5EScuLemx2rK7TUPdZ/Bq+Z2In1TBMo6xlGCqUb
n2a9+Qj8FAW00krrb/ZsePUMAP2Et3nWvpfVGI0cFD8lh7WmtbPmpSHbnmJYcjf/
x7j7U3PFvPInfEWVabzpT4OjOmDiw0agzvXGGZKVBVV1FJJsfaI66qpE89APWVGw
4B4TtNiBCoS2t0qSbPQ/3OPbNJ/0VfHxPmXL8Xoa9M5pgyvXxshwkESJ+OcEu4j5
S6jRLL1XDc9BVZ9nu4rMXXydCnCUJYjoGUd9M1Skr3aJeHK3NPtDJvo/LIkSW9ww
+oknfE3ORwPPL2IVwAIpAKsEjNhVASEw3tSV0OmUgM5Ts75Rl+KOu4dtsx81i1oH
w8c5sIoFJYEBoEP2OmKeLQCxs3L9+y72etnG4wHUKTwV6ER6LRbiwERTp7z9jWDP
ng9wP10LDelXmQX6GZjIU+v0MXT31nAvofxHibkWcytpxdDsPd/Xydau9AMQDtK5
aJqGNyxuKS6e2s1d0lBm4kE0S12rM5G4BGGhCCIg77tsHnVx4Wjdz6yZtn9QLs3r
ixGGpHSnrEp7Xvu2O+RO+NN2LaUkoIQm1dXE47+0irRvPsVGoL6o9mCGquHwmhAG
A5o9/pBC7wmT5pskfbCymjUbT0rNmRO7Sn6Fum08pkmF3kU03x+xMLFdiqDbm3jR
DmtuhqkTdYAaoGN3n7cfBmvOWsvOjThj4RKa0r4tfeQd5+0/IIw+IUat/zsoXeU4
k5mRaYAB4xKP2aVfKU7vHHSsQtidVPEC4aVGcqJNMBw2MInVvwz92ZknHikP+PP3
sbenaTpCSCdrNRtYO57VgvL5PeKiyZu7mr3wiff7XjDVYxAJcOebDdYqROk00cRw
d31ytWg3wZj36z/EOlFOR0sQdI8bV7rAwhJgej1OccBz02rm19Tf1oOrdU2QVPhK
SbtVT2s+pxpzBOd9U6d1gs/dbCH4/H11PPBcZ5/T2/6s14IeHIG1vOIo9ZAP/Ph6
+tqExst1B7WyFgaIPWJRx2fAei0UeB3kPemES36BH6jAUzg8hi+jWBDNmKkPtPZE
amXDaeUbVwpRxj8bZagzvlq1QWCJxzDtHFM3o3luLiTJ5J46SiWY3EXtepLuZPnX
j6kAmH82CnCTDOup4QCFA0Zq0elgA9cVY7gfMsvGeBeXae101UrW0SbETdD0u2a9
D/jxi5LT3pMh5ivsCncbKGZlA1XqQ/LKt8O9/g+40cwh7AfZ3Afr+03rj2ZxslQk
gEHfD+F33GBvATdZqpN0lXAx33yWrCcJPuyNJjtXzNBHSu6cKCiNel5TQCt3X56F
ODUzukbhC5qJwP2h8snJkNzRV4w8pIGmulVAGq4rH7IBGpy/wYjcIVqtQQzXqbPn
gGme2I/cj9mZsDHjuCVI2ioMQKdpa1Yl0oBHlfb3WOD7h+84ioTxMJGubLXKGClF
3UL+MpCzA8T/MHqwQqoqJ63FC5C8z7skU7gT5hFrsf9Sh115EBelfYk8jmhR1I9b
L/ofabpTZg91iYWHBLSDJ7KLywifbnn8+oHfODTGM2g4ejKvvEPb72VlJyOOm4HF
ctvVh/NZLlVAh8uwtMEbyUdbegawNqlDoFSdC9pVaW/3U0BP/YwQ9ymedHdpgmXd
RyDZZmukewoFxZ3FIyz9RffGM6fi8vnx7EFWKdgWDKNoRZUItpi44W3b9LonFlxq
wWmsPIYx7ZQ8IuQsY+i9J6XM8G1GTvkTpu6WmARxgbYAMR7dwh/wgz+oMni0URHY
r4bi/p+NKp/6cUarlzsV0i8cSRBDwJo3JwiheYMe1aCEkLUigqGsE6nvucbx4/Ex
9ahC1pPiy9EJlJMc38amOJ+MZFPIyEC06C34NiCVtHgltZHtfv8synH61+6GJ+HY
l9n8PWxpd8tYdCj2xDt34nut6Z+uUYqz0004USxbpc5MX70pAds4S0z+fBz9XXLG
ZXOm/UAJxG2W5l1pAmaXkwx9OVVztzNyjzmwhsq6h9YnalVRdfW/bFdTRY15v88r
KUvhLaG6Pc2Q7hAl+GF+I4RhOw8mbGfaH37MN2PiscYPmFG3u6TRHNtt0hzxjYDA
vx7/aY/ovXz9F6HlT5+UbK5XN3pVahZ276PuqYrAefSIN8iVMTgdAhx4F8oA3+xW
b/L/Zf+EPQChjIEn/he/qD5cXPMeXJ7dRHBua1ReI9F+2zBZlLIMIhUSR070qs7T
rOg+jJTwxtGA9rk6cCi0yAxN9hkY840QE4k/eFx1DBHi2e4ZYACjZSbyf2ecHMLC
DVM0E1jvBwMiseNrEGuRpLRoCGBPD36lE62xwGGcIyYGdsP+1QAcJpRUcnVJxCzj
rKqikF7+abgcwmnYeKtt62+4uAgsfAnOdpaTtCrZMyUzCoSHw01Ld9EPymCHg2H6
oiYmXpxKypt28LT51uYCdFAYGuRSzYTeApeNVmoZJO1l0k6XcLil+hO0xuwmHJDv
8Gbeq8gimohfq1zSQT26X7czKWrgsngcNoMcwV52X8/yPwxUsm1zeOUob2IZK8E8
iS+saQYdCM0TzXovwOoez1vgMmWmw6GaeTJNmKUpWI3Cv+WYM9sdtsBPcWYzw6am
5E41XiZ0zRpYUjE3eORz/r+crsqRHZetq829xkqQG+Vxls5U13KvUuEJnJMVR7i3
uby4OGnXUZI+rIZHwoBxi8ta5/pAX7204cAlyGZ58Tp9WzCscAWZHYBXCvSGKDPo
JKWNBX9nSj35r9rIHPv/kD77mxkbbYBX8EZAOcvoJ+LmrU8Ho6Ev/ThwzdWTm2v0
OL0byvk8kgi/Wqs0lkJoGMaEizCnl4zGXmbk1y3g9v9qARhfRcpwviFDzgBQvbuc
8Z4LrDad4MCyrXqx31cudHVCkll0ZMluK5mBgtZQbWr0+6tGLipgQh/1DWOjdFzg
9UwejU5PVDdE2eRr0YYlWSPY2pfNTR/CirqjSBIWn+JchhLblpvKN9S/2gXii4jp
qy07g7RHubBynocJD3+V9vCyicvXjdK4onUNFCWBSyZbbcpq8yn779EwPeFoKfT2
bZ5eSkdVW+OPDhkCGv3Rw9AhqOWcuoetihkebTbxE9pEhTyuBOqS/SmzDT/MO5LX
e7Y6RVapu4A0A8kU9/eE1Aqq0KUAJ5bF4cjK5ST2x/CP05Jyoas5oGSEZpQQIIVu
NekV9TAhQaBj5cxhM4r6PCkAWpAEUqW2vNSXQ4p1UjgbYjBh9ElIxG6FdB//tNVP
8L9bxADT1xtjfoD90/u0dSNeS+/l0JV6aqjvCLzsoDz5xrZf6uGDSaeKza8tquSo
WR6Px23tcl82WTC5IhLBfnoJMqQDQTW+Y8cn4xccu8sCOrxgCf11Fo/RX+9Tp6oS
sasT8LRNuAIFP/AvngPbvE+oL3wN0HeOdvv8VNJn9b/k3R2ZeomcsfCuKYg/JZpO
OVCum7lrc/l3m+bQTi2o0yJ8FFJPmBMZ/UD6nVof9fzD31p3dXewLqg/XcsphA55
pxp2Nikz5HirC6oe6gaizfGuu79dUE2+MUODsH0zCtHNfu+c18Mheh6s7RfP3tjO
1OAfr2dvLZAbBCSdCBE15wZ1qrlpbzE+/w+PhROModJyB7q1Fy8CdpWYbZsAH5yO
eFf8Uq1wrWzVOr7XCBzih4NvjbSSa/om6SKZgqZvfcG0S+D6TR7tgSptg5A/IoGT
uv+xcSDWueRlTMs/H9D25ItxzgQ2lNpGA5n6DcXJIcih1j6vtp+5+sjgoHag5to3
56KzvwvUH00DPLps4ven10ZUg0ocD3eIGV4HNb0Yg05t9cc0QaVjcmiznkDB/C32
k2cOOJgwX5xJVnC+Oo96saAPyUFQodb5mTefgD0R9KQ8XEua1idf9xgCb8oBQbxU
FmvuQm5kOlwtiMkgfOTw5aT6WYn2EdY/g/OdfJSIF3h5iZzGjPRR7gtEsMGV7YVy
MhjN2ovtk1DKB7fLPDSZxG84vyKiTMJx1skdH6oOIoKx4Py8unceCwPcciDaepOS
DUR8Wn10TdpiPjbLHR5x7T92RyIcCyDfNynSW5CplHSKY8Rq1QCacf8ENDcj2RzV
bmBxxXrYPAEQXTaSEJMtUvoBscmwfmNhtwPy9anQb59ri31B7AxiJ3uaYXJ+Pokk
wu86TxNIbQTKQl1G2vFe2jrXWDiQdxz7UQKhD3WF89c7itsCANFAth5U++rZ88iB
ck3RcC7pQv+6O+cSG6IuezT8BkBn+ZCKYWKAum0+/Q6DNYF3qf7kyUFrTGjfPfbT
ccqh7txYKzIAaQPj0kAo0S8UixBK57pXWmlFTvoCfBlLrHB2ZFbfYe+I8HVupw/k
gT+eZSSoStGqhk4sanZGHfBu0cTY8TGJxYXMYLbHogO8bgVTlBcHb9c/fuTzW3tm
V/T2j+4rtIFXD2qbFLaSYPIzF41tCREH+HogpvWGj+P9JzVk4gMItzvNy75sVAS9
QVKpSnopShZsEPwakK+1CeiNWRkOGTWTIAViruR2FjpttZfcRdnGIFoigAeXCNoi
m3CFMC86RvxILk07V2twtbtfHsIx1x/JigVZ+3kw9TtD4VU8LNnjQYz+qMSvUjSJ
VwXW2rDithJ6WOzCLMjT6eMJ75rVaqBYyTob86282EEqBna8JrtOgotf2hYJmG0c
t6Lqi1stgr8qAs62Yq+ImpNNjto1upWJanq4B9YYBZheofZhTthXLtupkT/fy/3G
gZcTgunJn13YPEdXXX1sIwb+0xmh0wfLvGwmOOBE7ZdCQYfU39quh2skTxBSqX9j
72jfMt3r5rDVoPb+B9wGY3B068FufvWBTx1nQl43MwkaKfE4knRHnQUDXtUQzJW1
lboXFXMBZRXZA33qXNn7UqCwDvL0XXb0ZO5jJGBBX0Jnn6IO/xDyvKw0sJVmUTF4
Jr1X1tTkzlhGvhkqijxGEs9t2Z8WjZ0XdT+pnaSNv3kqQSuzurUZhYI4WI1Z5NSs
gCjWVWf7Yn8vFfTIfQP2PUE/ZtwW+IvFxro43YfPf58/QV9QnUNY0z0aOrc5vXdz
Ptcrgs6FlctvRJdzp1HRmJHSedh92tDkJFBqHcSlYZwdxq8UkUuNFRCR5qOZ9xeJ
QTGIoB9sBs+geGxSIxjC77EtZUq2d6D1P0CwXVNwgosGPhnEXiwaoywg6lZKM/vR
WNWwTxVdpS8SXiTInft0N2MSMqsenPev/pTwdH8e1gO533aGoNFY29aPQXZdiLUg
L8mNbcBTNTCE5LGoE2x4D0cg3UdtqwqM3eiQY7sBgEN8lPyGtGzlU4xlkDyFQ1kS
vh9MKW8e2Joawz/oQUoW2kXPTARmzsPLwtOUGPyP58AWe2hKR7/e+7HA9UFZTH6R
NipCq1uKcEZfBkDnPrJmGI8EFX7+RCeOP85J1lEJM9kXpOxHyz7H+C5IMK6SQWNK
8O3d09Uc+h0fxMlTpSoJic/LfsV1wF9iPOnp1V37/usK8EHmu/KKKN4PthbFJRc6
vLC+uvskE/Wz6pexzLkPimypJTb29SpfEMaV/msPxk4r3quqAPmIB6JayXPIfYcr
SfXHgfr5r7xJ/PG+yggbpVgbp63SXR+sXqtJ5+zlV605YW0dgXakRNBwFfa8xs8b
mTR3y1NcTPYaI+ICPyWqpbpSPY8UxLFTHRryM8x1hZi6yuISs642JQ48CuXXAAeX
N8mJ8igF1xrTe1bZRjxOjrphrDRcbWwGl8fZJbrjXTLQZl4WkP9/0FsXCZujGRjD
DHPYQv0t08XEMWvU8zKm029JPOOMllYkpxJqmsQAqvuqO2SAzcg/0jLFkn/jGfkc
NJz8MYZazQZ01zIDH/t7trJdDaYs6gibOeg7ifFErMvK8PO48e+97QHqH+yuBh0H
kpSrTQHAOyKnwlsfJgrCZwsca4q2Yc3IOejiHb6fpAkYKGjhEoaU2nalgmGbfke8
Lk4KXHHKldNCL++iNwGz1zE27xbfMIIdb0a59vRIRg3bptwGQD6RdR8ZG14ZXVod
kocK+oopx5V385h1gveP7hvMIa4bec2rE+kv+qGALIiiiI7tWVXwqbUCumXgfYvA
To3K/ETfz+MxIMwWRBydwE142uUOyr3aThZu08t2ZlHTUeLGmJijRhEho0b1sDgi
b/FoIPntXBI9cTMvkTxubU2v2iCUeAIEBrhdB//2DOYA8mV4IfxahVyIEcgNbNpT
SZWnnFBFxO2QimqArN52zimVp4eP01aSqbHoCmVbxZQGAVb9gzOnPgirZ56N3/gl
z68lMKb+pwGT93PUgu+gmimYBOlvqsksohgTmBE5hL+DKsmvicYanczf5kieKmR+
jWTBJTTp2mhyMWEVbB22u2RLv5pkJaUC8vl1+9w1QOznG3cJGKXqxpSJXSkXc/8T
vZcWzLExjqAveqeGUtT0T6+5lFJ5RAzjYt0ECoe/I3/1nSoR1hwIsOQrqdTHkMJC
Wc21oprPaminFnife80FjdgPKa18rSa0RgAhzul7Os/19WdK9kodVkt+Y4ZnOyxL
y8rKwiPATtjh2/I6RxHjxdSi2UccflEOr9y4jI9A/8sxYmT2/LkFyEvr1B9NLqu7
sCKzSN5KO4ILAeID6YJkUEXYRYViMyugkrI2d9FqXYVZlM1BT3Vrd3vZ/4TvN2Ik
7i4+ZLO+MF+gUHX/GaanWwr5NAPB7pS7k0ZPGd+XbgVkTubloiiTIbjkhB6hyLJE
42O5C4ISU2S6GpWQcJCnR4MaAoh2UqAT0zUFY+Mhd0i/Kxd7KvJkkDcYZfE+bs7m
wkqmwX4Gno4DskDALlQTDRyMNeb9Hj6lOqyCUzIELKvLIVo5IpIZ3e9K0OTeos0d
WXf11y0RqNOXcvhrpoMseo+EkG5mnBgxTEeHWwMrk1f0EIKiagLYVjV5nAez8dWi
ldBCtnXJVlgfhtqQ/zmKaiv28M/kGIt0mry4w7KoCMCqFUB5MB37n4Cu48bAqd2T
7tmwHXYRfsVeiDQNTru3BNwfxbp4d5/lKYgvGo4vZbbTsme1bGPM1Y9V0WBBuX04
2/fHTedOYY++Vio752CvTiRE0sOa4JKNyZNq5h8MIEq1ya/2cCgndt1ek9kNJsTM
0FNHODBrgXPaO4sSHOYazS5BWM7AhuAvnLeqE/bsbC7gj33oN3E0/kZGVgvXPxv5
HhMfCQDdbu39X949cp6IDyDYDj1fwONsO484ffJIKoBMfi3irQLzYqamex3a1CNM
7IF7iSv/NYDmOEpmRbmJcafmMqtIPlL8GZx/QVgOGuT6RkZA9eoPCvYGhzawJXH5
Xp/J8GUHqHLudR201eotIpct6/d1gXe+XYB3dOVUf3MwE92Ou6ORsgKGEKh6bW4j
OurE8a9FWSiJ9h9CMEWYK6pQLwkLNjWByJHLwS/GkZUF3OzJp7NcYuixifj8wGsA
9E6lLFWtHg4YGBp8fbrHFG12BIU7wIv71UdXsF4hNJja7teix9KGyhRvveXrfqSL
kDm/Omz+xef+Qp9xBnv1Px6QPljhO2pUmDTAEYXS8Q2YnYqf6e6r67P2wVnpifNG
O0bjeV1EtUwJ1u3Gtx1CjJ8aw6tQaPGuNsNGOrV3x1LD5Cb1WrkIdO2vFYMRR6sv
hcHBSgZk4MIJuLYPobGxRH6MJkRPG33CU3vPxmmoTp5RMkNzGXZ7y7x8XZAC1Qj7
L48/8uaqCXUOq9qI3+ypna89mdHgcQ0mYiG69/jYuG8wzZ/u4mccHP/TvPsqOgB+
ynYOVMf51JfviuD9014gHSkKV6I+xkwmwwgswv51StLA7KQh8CB/CVGDcLUL9LEi
1AKSpK5v0WgM7qEslA9pjGN1KhjEK5iU0za2i7cj5I3wQiLHyCW2eFH5CgwzZjfY
EK9U/fQmlOE5zaFgeSNk336CIi6l5yEq5n69sG27XM+ZSxDA+GgWxtsSkIbyr/Cz
zb32vnCnQl3kp/Q2Try7HmhOHwOQ2c2W284tkld8ZM0PBXn/krPs0axqHhYapqzM
FyrETqW+d3YKfEatlZN53BarbBIpl7uKpJb/QXT+nEkGtDOkS+zdMeNcCvuIgvaf
Vu/MuP0cpX5ne7OETYvPYoAkbqP7pKKyMOUvWcDdEV1YkSL3uHVqPEW+1Ul7DFTe
nrrirtPo3+RFVYPY80qq2EHHtPVyHigL5AW4JjxNchYBTd0aXxeFaYmuRsZzHF3O
MrextB5b6aQOzErhKuoLaLITREJ12LkNYFwfNW2R+W9dVK8d/gt1pvceT41Uuv7O
JhDXTOnN26bbyaXfeHBXvHVIT6Zm1MaQAa99vTnSiEpjiE7agyYxBnbgP0+FKxFq
671km0uEHidRjxQFyIjCVo2+OAnJeoDFCEBbqAVhOwXA8BHcYC3shEhvcJhs+kWW
gnBee4pQUN9FoPTVLivb8z4WaDFprTgKjronHWVkNoKe3hoGB+v3k4uPBd3yRxrL
p5+GmCC0080LuJyq+hFVlfqtlZxs4K8F/kaZDvhuqEK6AGMdnGaSHK9/SWJ5Cr1U
H9OXtzyltwBw9+z+xQUd9l7tDsyGvvwstp2PYF7pgBVsaFk+pKmgvK27LnqoIeQL
ZtibZ76vxa8lAO83/x8WaMt2Ei5/3fCXngT30LMReTqFYDr0JpMkqrtSi6NhXKah
xkJSXAOyWfTiQAWIWI5Y2IASbslj2UvJuy7Anc24SqaLPd7NmTA8weY2UxpBqu2M
soFPlugDDg/vdqssDGDKdj9TX0yIKFUnIIsqDTRXcPBIPjj6KCBp4mum2k1kVOpZ
UmqxHWh5WQ6JcswdyFVPpfKchnXgqFyIPlzDV+2tiFNAfjyJS7A03GRQpQTKZKkl
nluoJPsCjBjDP5kyq7N2pR0+QbOrYRXMhv/kYrXHOghQVtGC4H7TUaMbPxkXO0gc
fV8DyESf7jXN9L47lK52RsDUqIm663a9GnmrlOohzCggQq3VS4xc4021b8qwa6C9
SpjkT5py1/g00JORc+8XJDyn7sCKfxzfdEaNiPLGnd1Eb0jG03eNJTs/vsKUIgKO
0zoEqEMe3w8zLYi8lTEKMzYeqT4fRtMcu97qbKIwbDrcwR8+oZRYuoEQJvAQBlDb
XBYk5JMYo3iCqGpWcp9FTFVimtGhUgc2U+uzD7LoHneITPlHaMq/kbkmLqdQJCWq
Il8F85F7U+UFB0xgP8Zicqd2ehQGQ/o0rfA203meyDwu1b48a5DTP4Lcj+tEecX0
CmwfXdQP24olDmb6OVDJK2FlVpHMqZPprb+kC2tEdEb+9YG7OUh3Edv5hxs73qlR
wf6dFLVIa4YDVTkAbgDAIanEmAfh3mc1RiH7mx6Z1wXwuKMaXITB/07gQ813chEg
ykBum4fzB5L5XQFt+UExDKegDKhIeXlqetzYeSwiSq8VI3VNdYMzmYgfSi7EJo4g
+iJ36wwZA/lDcecOwAQAWJmHAvDYUXW88lx4XphCzjilfk7uoucSLgi3OdanrRMh
GkI+q3Z8UWLb54Xke1uya9WT783fy5OyfozZgh9pRJldXhq+BJabpOSz3j/0hxVk
A9taoXk41wQqs66cQUiTfn2Qdn2yAl/qnokMyYJfSRFzimKBeuDooLHouZw5gnNq
Ky9LTHWvOSb5nZ3sn8clrDVxYxvQsr7wEN1WdekfRS0zHIG1w+1vg+MxwDutOkcK
zBbud7Y7W4uJCqFEfQNvhpOHdoXCQqzQocc1bi6SDeAPtDIdooZF6RvBP55O6jyv
OMdB4daSrDi9f7M/vuIO84TQKx5hXQsrg9DeTtTTFhbTiY79zaOhYQhdd724bfd5
v2NnKP33fuqdvxgGa5pypsyMzdLrdzo94t6kIOybvOMDpPvL3+nCLj+1e6xfVbl+
7DV/ocYbpPq4ETDePdILvoeQ4Y6sr7ezq6gZN6+XbKPjm1uQMtiHejEe7tI9FWuE
sIhy/lg39spItJK57jgybJpm5DqW7s01Vs2iRGthm15SLSz/opLgm7Rmu58Yxn9W
9kS+lxJOuYjfMDwc/glRIqhTVand6AthobWBNaVJdSUhebgH5RdBMP2tk+aooBWO
Ohb8FiNbtW/wjb1F72xgbWLfpcDAOrmWGSi4B/JVHLFntXSfgkYanCHa+S/F1qIK
clB0tzr/jiwWY8eXb0LlbL1H1Y+3AF+W49whXk95I0SVYzbr3XWQ6pWVEsP3E/4W
O/RI5pjS0f2tUVLYCbfnfeAsdVSXxeVa3W6fOTvoSzkaGNHN+3MqxFOrcOuH9Lec
ZSAoo2uwbfsRunQEYZvRkm9eD5EEYgTiYunRjM7Mb/DDl4zbowMK8GaqcjwEeOQx
pn27Q+M+6Cj4KR9x6k2QkHpfyugxtX43AJr+lkk5m29m6nNl39Xk4gRHyTp+mnL9
nE/I/0mj9RcsGNEDKK4St8cVajojnnpP+wtAHFnsjF+Fwu4EKmEEeOkhmLQxYdnS
jXAiwPlW0oYQoDoscqJrqR+nnYCt7Ugct90ZArN47dzbpM0IYcqN/cGHa/rW0N0E
dhz1i13nhLcHzlTHlyT3BS+XoJiDagDowCJ61OwqtAH8B7tFiqr6e9K6goPw7UhX
5UWCR1p/efI2TbM5uzmygKb5Fa3B+B2A8sskMr+1exNVX+Bvb06NzerA515qe8Gi
MFjHwg4H93/oVy7di1AV99jN3Adej4WLIZV8tNJTFnFD8R3PQ6t1vVfMkvtgeMG3
bhwR3AaAIsJGzVcN9nMGMdgLFW8WZE4/X2XVVWq0baDDogeg0j3FWg9dRLqi2my9
tR8zmq8/c6UiT/XZu9n/AYaG/WOfUKnHIwhSy1piForh1l3u1yU2uLCBpv0+SzVi
o9AMn1v4vNmjwsstI/aIh5UwDrWPV2v9LyXzCvvePim8w+tVNGfenUyzMmKqNc9j
xSuCILgh3bS+tovYA/DMZ+/P/p3NfZ59KV4lfwErA/WfxKfFCPDky0uxjKlATt+N
ICi37T7Qeam57qTchuIS75lnJ8pcv6l2Ft+ViNK0vOroGqlydbTOTZ7zztkLLIHA
XDtdDVS+wSExUuYHK6bKrikqTgfqbdpYA079FMQWX5frx4R8rfHPvo2/rtNogo3F
Kjqa3bqkj29ZAk49FJst8Q1LbTQuWdCJHNuX6Jh7UZXlnf7IOTMIvK+12ZacuhhM
dN5NQF61E+zmvWN8x3ACQ+G6euTD6rAb8WGeWqt+d46gLIxVquZuaryfFTwmw+WN
qLL6zCgSBqsuwggmxmnnjCvL1IEP+8xGF2K1j58TD7Yv2oBD61oesTYslXLEgQnE
rx453GLBFsglyaQLwppPZjsYdKBxZg7D/yqwoucTLsVQCjZNbVvGBFkm6VZbDzUO
gViTykpq7fQCzI2GHDb8FHeab5poqc3TUVL5s1KYZrlCsvIriZQm6Pd3+YzaTsbM
RWNUeHXLWh+Q/VukUzmeoMj/CoFICD5a2vXgo5dPkkAZbEIBIUS0n97OD3b1ks+T
v1pY6jajn9tdiyOUhValeSk/LXIyo9sqhDTF4BxsJFIfgC6TiMILhhcpiAvQz4bW
lMC7w1y0lrH7j3qOre4uDBAzktOFHReRxgsqXxAWsSkb0MaE8UJJfhmJlNDK1CRn
6SUl2RGhis88WaEtCYthZlaQEdga9i3kY8Z/lfzik7TXLjDtUHXWtacSt4bs73oB
bH/V9Qf5teASiC7Odkcj+sOxy6DTbFRKbD13kBPRFhlXZS4BATEfDAdOr/UpvcYx
Abl0/JU7Du/phWkvvIzN4w3unnTRF8135xxvG/skl/wNg3KW0UWOcM8dvfr1J00V
NCnprDLY3JD2bHsTqVMdk87PfJikPhIF7pBHMk2G0rTDW7+zodiOS3jzr/VnWD8O
B6yHoIzghqx8LhfG8tVRzJdDxuvnyHnebtmMCCmWaCpZXRp56cAVCceOVHDS8Ycq
zNMcmXqaXFJjtV6lcPYgB86vzcjSHBp6KK1SRPBmLbCjfGtJf2UOWpBH8GRRtgv9
lWl/gn9PPeNnktzZkJ32Krs3swQIb33loH3t7z9/WSED3/+UxXlgcXiuBPazzC4P
0dQEn0Wg8wxgcdHDTq52bPVfl6973qKcw4ajy6aB/dc2/iJhO/50E3C+guePU7mZ
B/1Svswhcjcq3DO5FzYKRF2Kevun9VZf8h3gTqVHxsYc5XY7psa8Bb5PSbPPNa0B
AY0kuv7qKSfQhuQA/F0b5eS//RX0otDKFxSDYH+kac4uUYfsPTUu0bGsOLr+zI/3
ddFb/IG+a6jEyDIVmLvtJfHgQvUuaF0FaYlXpj850y0dBIZSbS8RjJm3B+6l7PAt
/XIdBEGsfli/i3fQt69/ENVlMCxDROZTxAd9O98/HxsPRcB2Jmk6DayWukir0QL/
K+6yK4LXaRao0lTcrClhAEuYE2zu33t9D5dhrc90VgWc7orhwLDljfxsy/y9RYt0
mhaVwhb0gBroROsx1TuihxfyCv5YBOAKN3MZEfAB8F0/JlRzQOxlZ1L7hPFrXHGj
EoHBAg7iOIN15ZWcfDfzs79c+9TYFG9EIRhQN7mvtcuYAZYGmZh4P46IUsEnEmUR
uIBVnEJ5j0ylhz3GLIlXNK68edUA6pzHpw0GvGSp/juxcDAoSWOmBuX9wieD2krJ
S0PgR/S33XOqPY1zuIttn7pdh5z6P5QGyYhifl2sqoshc6ZNX0V/Bv4r0iAKDtpV
KC1Nkt4ePUQ1NPzroCHoLsxFjcIcpys6WOpr+Xg6d/in6Nqwjc4wRKDwaUDuS1iD
EsG+NkYeXZin0N7VXgbrR/ndlsQ2mlWHnQbGjBY0wZpnCXZzA4aZLKEMWx9l8Kfa
bCPycu35tfGjfuvt8wXeGxN+e1WXdZ6ohLvJi+Cp61ujxdpOHcC2SqaWLOFUV2BG
ss+QBpHT7bHAWYLJhrALOyMAoDW6YKNKav6ECDn87IQUKl3KNeWH8/a1sUOCusp4
J7FqpCRbTGIbDQplVE3R9h6jKcIVhCqj2Dnf/8XFxm5kHhJI5N6ndm5QGohxCjnp
ezWOz69Swx1grGHoGs8fuxFI3xLTGS1ZSy7ln3Uj5vnYdAh7hZlWT3Gz2e8v2tFz
/MQ8sSu1+U87+SyAodNo8NtuKi+tioLasc9tPb69JhLLKNty5Tw2f8xjREFBJ44e
YSNoZW21792L/KkxzCFIruQup/k+03P7WTBcm4D2Nyr0JlcWtSbWCliRLkKYoObg
9MbPcUI3x9dMgdBI0HHe2cfi6V5KfRFyXopX7Bcq9u289fgsiNyfYlwkWWWHADV1
W0E1GWV3QxjqvII0B7X2m8VTBU9erggZcwuHwiaY1yQ7dnIwTbcYRi92Ic26ZBPs
Rp4K1zb7amk/5L3s8sGf952SytSyamaB/fR5kkJId8ISeGIGh8Cmnh05xdC6LA+x
jFn8nhKFhn5TOvxMhq0BOJUvXj6B1QzpXE9YSwx55OAjMrX7Kf2EshGnLNJoRZ13
CVSFD830filUxVmvljF4rbDJRgXiqPLQtmz8dAWBAjMbyyqMRomAGFHEFp/AU2gm
BwKGooSc3d0bkQXTl1oJUtFf7At7548JBj2I/4W9Kad+PZIq7xYpI0DUn+ARSN4g
enmmvtdNQPGwz2vXsjUNlok3yv9PsSzRDEDBmMpEHKY5OdBQ8dE7N8GThKGU+poD
Q50f9/xgzVUdNMSi6Ck1wHEMt6d2CitVWZUB9/tgRQPZxWrHsttGDcFfOBiL2CHP
7IY8rGA4T0f/oIrAMrmIDN4VEr/APutburfZVh5guCDdZkDAkfMohgB2HTaFIdtE
QWN+3dZ0IMDG3t8lsrYePfSCx1qXRm1NDUG+UpWWA9X0oN6rGcOoTZpnEK6FTARD
vbqkwFnqaV9nf+cRODhe+qUg0+wZsg9AzDRzyzS1TvB7UJSGHH/X7RbgBBY0HKW3
jNedSLeBTjesi482TiQRLPG2BLYdCcOhCmRLZ8ar/1cddGjhkH7dxNpyniD14Ndm
zvNl9GTe0wMuCDXJqXFqZBaPynevnA0Ke+wgP9YA+W0jy+hKEVeDTEsyFFw1Hqml
5enQVPkWm6/r3B6gZm89EK5otslV3nZa0Yv3N5Xb7NHAk+7ePfO/M60vT5/k9YZe
qMEsYdbTXxqHdSvbl64oEUYYSZBERtSsygnukSXKE1HWP9iTzOWBC/dve11k1CGu
OkIvWH87XpqCTsQTCTOJ0n7fq61i9Fw8KRmY0nBMl3HlmhyeJ37llRWTHrTN89Dk
wwGdJnROqGAUzmE+/8CXuNb7zBkxNRfWyGFUQpV75wYmWo0Zn69cm71pN5h26lR5
sQFKt04B2iuk4dEKsLovWdauejFYPwOoB9f4Vlc90IK3RIm58zKZw4I0YA7HGZMV
3sY2W15b3HY/qJ7E23QpgzfmWNHQeb14RG6DrTZPIJprUwPzAps/RTWJhbSBplMo
X4xmlrNFycfHNo9t65vBiQ3vkyQYkWdbR5FJoygDagsbpxkzEknHO9c2rbG7oDMj
6FWoSqT0MzCsbO00vCo+QrO3qltQYyaql9Idfqvts9Y0wpTGZ/thbSBRXMroR95t
t3BI1RVQU7QoPCPbD6LeBo+M34ljP552uKAZrDBVWriHMlVWuYG1iRD6/VOsSB+x
OraB103ZiMuqtv7OQoLm92qLU9V6O+VE9A0HQPPd5GfqAr3YXSVAvYsJd/JPwV4+
E+ApCdAuqr81SRdA5BGBBsMrePsw3x5mFre/nbh39n3TdVIwta3Ox4O+ckaswTo9
8McDOeIombVM9anL3d8JaMkIsVfhUb0YWOseWkTYzY1r/1TEnLyYxwsIQl92N0q2
p9g49hcaDUdkJ+8UQQih8Q8AEuuRiFTz2bcBZQ4FFMStiMtyaGXsOtK5Bf7GnZ4k
TFM/lM272so0DmT/9yyzi6Kin56B5+qgeqdU2lobILMjHP5iiudqFH1ms2suBF8N
eACzghJF1bCXsn0G+axL1jIRaX7BIPX+SfrcstAKHfV6PzaI4ySMVwO1WoLpfLni
wknuQiOVgJzS9s1oZIsTkkl8Iv8+qfFMK7WZQvXaUSduQjDHZhj/DiNXslnobZ5L
1CTZ16CnRlLzwet9Fhni1fq9av0uPLvAvF7yiMa3B5zY9lOfVUbvwmxXhdQmgBJH
joOjm/ll0n1p5uMcNUmIQJcKQpwkY/m8kJh0Ivnsb744l9N+pYVqae+zRm6aZh2+
xj82p7JcoLimDEAZfl7ZWzVEifVWb7mZkZfw62s84E+J+J5iY8Un5AZbCpRhPbuh
J9jBOsGT8YiDwKaqIYfcGgX+vtWftS1HNHGJzgSnTAsjJrVA33bK7YNtIn/q1C+L
7T+5x6BbgGUA1qOxue9DM3wDtMrvEsz2d5yREajQzp+eDoN5oDhllDQNICNCeN4s
bNPgUAxkuEDAHe3CHhPx/DrGcWbLbSEUpxkuFW8zGXuGS3cPssZH+H+IrIYwHyZO
Xbg5pov2lxNgvz3eaIYMiqO2BKsTCoZiIGVKMMQ8un/vJkc9ZeQgl2/F8gwDT66i
Jn0aiAWjMa29JR6siL9QS3CMR6oOrpEz4DlfoWV/od6Aq3ljBSGhBEfBTeq5mHCS
HtAl2NM3WGkQzq4jKWatvDNhHvG3i5CDFEYP8n8C6Zcn79MPjmLqm9lFreH9DhyU
0x9huk1UYcTCC0yiudGPeubdfdmOYbotmBenXWIdhvQChXvYiQ5Qvlngu2i9FXyO
naP7RxEW0bOmD5jX1rDaHCImG+LOLUUycVm/GsRXVMGOK+zs7sz0QcOlWjc9bHF0
RsmvA/WgIE7mWKR+hiJ7ON25KS8XIMLpKG7/aWUWDqMyT8NIlMRxaO0UKMTBR/69
Ws1jLcxxawanOJan+RqZkNmXXOWYq7toCjyAJIPUNGhMthRs6/vF/hWM0E2mxsr3
6FFwJC/k2qMwOZgxm++WFIhaD2FXwmBTsz//LE2gcc+870CfU2Mmyz8jRwQOHB91
sVuTL1ig4b0XqO+7G/mUlI3uHoAmUDCsXBS6mrXU7r7MjTL5j6+jCK0WhC6gx59P
qKyTt02/YPEvRYk9cXSWA9WR3lFXQIuiYaXUyl//bsguOulcQnpatAyDVGGf/LvV
NrjYojSjCBMOFFlCqMuPRhDepBiprt7pnmq41FTLQPwlvhHUn0mtgc+5zyJ1OxrA
dbbvNmQT/WAcQ2ssrJNUDXLloZLtGUUw6uAbYrH42gK+oce74Kfcsk8Z8vH2oRF3
DBQeh/SsBWCb3ohcGohbi/crk0XrAmpWiQqKKzCjUcEIzADYabSVNvi2akYU6lTD
qCdS0J5UjJG1+dsFQsSx60uWFez1dxvpdllq8Xs29TJwtDQg/y898H1pnbroGuvL
6sBpULbhZfSjge8o+4kaAZgncM5FeWyooi25LVLJbn3C0tV69Fe0JnupNCyUIfJU
aJoVA6NBgVsGaGVVJ5gg0DkYZqb40Rt1C4DxT9yT5twDtm9KYt9CyaefEYVbVJmK
cyl7myqxoGXY4E2V5j/k21N3Cmwety4mxi/Qau6xc2P8bJRkn1awgQZ+vEc5HD1s
6eBaPD9bQnoERUb2jCbMXfs80yXmEEa8eeK/mmWZg+uMbDyV0i4Vla3RT/Tg1Z9i
LbodFIRlo3+P4pTzR0H80UVb8Z1qaVpDXBOIvgl3AYlbeCR9yfrEE3RsdawKDm4e
ibOU+zuZ/bE9Swvqu8/+mANKO1NwRRPzCsmhpgOJYHexAY7Lbd6BaZq5UYf9HXgw
1SQ/VMMkUFNx6EKsgei9KXih8txfLfkbsqrrrcrGNeE1asOHGTsnfELRBt5CtJPy
KFQOQy/7BIA2Fq323u3t3uCXZekf6z+muGg56b0FcwFdZx/UuLVvmaLEW5D0x4TM
JUWg+CHON2nyS+s2l4+EnmbYqkWBQfzYXbw9SIvcAkyPbNedRLOYMFOXG5QasV2g
+pYTOIOgDOgtlgPKyReOM26GYax87TabapR8L+CznA3c8p5E/e8hf+dHXCUiwUAK
1nIAv/6wDLqG9ASZitX8tlsY0IRq7n71sx4Rv5WVMuUjzTCyv44aQbJIX+L/xPqG
Zn+19ZFVon6sDfwGYc4lC5915p+1b2oc8f2tPkEbySpLzN8P9nDrKaR9whvCj4ox
ZdtnJ+93DhjN410VkzgNE3puOeIg5iq8vXOYCU6RfYXyi0y0F5Cbs26OcCBSHp7E
K7LVkV1VI/O6rsqeASk7/GTDa66wr78nQmiN0GoqE1xoFLZ6kmMtO+wa6Bxa9vcU
afE2q/TVReqCNp8DQycekBwpUIz7MUs6BQkH3AniEM5zv4W0FIduZbL5HreofMTu
8tCpbffXlW5cUPE/wWa9p9rcoJHpK19Wf+q8UsZfCKopbCrf/o5zCO4myTjNvPhO
Q8oHvIIGV3Suj/6E8pvOlbWGnQd/JBbyqMV4j/oVVAMq6FiNIE5l9LqZCKXKMJ4j
3wHCd0txDZpnZe7nbSlSVZL8NTFUgsMBDkc2s/ydSEZDHHHFy2vJhsclOQlmkq28
pJbVubH+Bb13t3/Fjd2zn6Q5ptuRjpOu+zOFcsiqviqW3OduISGX6BwSXUKKRZPE
cxahgBkL7jWJvjEAQKcPH+x6M+WPq16YiQrk2MMahJiybhw7CKmRHf94s8V6bICD
hKf3/Om0EKHTPgYmGbN/tLmqM6q+QSob53OmbGCegHjfdZFZ6PvYMV4u08xjSPsu
PXmcIz3kwYvVfPWTuG6RqFNPXG1zxCM88NPopBUphe8MJU76ta0Gi64xk1ozyB/y
AZXgKQphJyu/PcOij1BQvleqxh5CN+4BSyul656I27V/sGghCADDS/EzAaXx0hMU
yG+kw2xA2RD6Yr1zQ1ZIOUGimagjnDbNpPTwbwbg60mOvSYgdSd8nn79Au5Z5/Cv
5QJ0ExcAAf1wCDsppgIFxaT4DWaxWiFEXWnaXYf8vv4zjkxH2scTsziVy0gVMkUC
4+YnKOpBEdPbCqh2pF9upeBigMfe5w9D9g8Lxlzb19p3Q9c7XUREPr6RH++rBUSJ
AlcFYQuAtMouNtfaed+QEjgwDAZX4B5gXemgNzN8S5nze/NP0IeGGMnsbOQPJ4hf
McYHAs+54HAdtTEBKFbjB3Bn4m9SlKwGcjVIllCRlDPA/0fZaUZGxKC7XbcfNw/M
/jZhIK3uedSIeZveZGAXYmZadmXmNCr9kKPypzd6jgBemRyaglGqVCu3Qh+13jPY
mEsQFKa1DswAzm5Mnf5M3UpTK70k222ofFAbHytZ3sDJ/KGeOed9NYKnWxQwbMtc
hG7V3hVFAt2xoFlsW0rFfhcABRfQFABE0V7Td2UhEpuBqD/O55+VEdv+xl1whaqs
Zz5EhN6UWsAmXJnF9CuCZknHnRWAT0Hv4xcLUt2/UY54ubSjkvuPudYW8318B5Qv
YJQVZ4VdmHDa+Xpn7xpOoKYzjknaiitq1TRado3BJQJg61iqAQwUna/ttKBJOat2
6oOD2S5rvmpV4YzKWQlbEQOXX15AFOYLvdMqZ1588hKMgA3ASSgzPNTd3Bn3udh/
ej5WnsA6vMPU8uVwih4jQWNUjy00zkOayF2EfzW+67C/yox3o1DZvahE2jkxpFhH
i2+0yQpzQIrcpOBYsOaLL096P24XUVa3GGsO9ajOJM+0mgY9dK8KDJsXwOekQBfp
KSovhbEhOde2AXe77rtoEkc58a448PdJSc621XoxrT73osPKJt+dqXkntcvd1lcx
qeQAPW6KexzwIRaclod+pYZb9FUfzwlGnZ8XPwsubYj3rvsfHv7PT0oSbltzXIFo
UpVZxoI4d1CGQdPmz31ZI8vjTZ2Gop4LsojAwVuaWHTfbVfujIkOSe7ar0qXZ+t6
W5L6vVXpkR8EU8YMI6NxkSyglHuwZbATFTwrPuBzQSDcxibq5xAAcxjAf6X/LnFa
vWaq0rJbn+X2qDXjxETonnnzRLafbk9hDf2wqmv0MeHUXjv20+VhMsEbIvZps3Xx
iMxOFgl6J1L8BSnB3gIEWrJNBxTQ234FItthGzfuO3fOFia8x1g9vN8IJ0MqePS2
vAVP0VaEKz4l+paHB8kfLtn/iXlWd5uMajqAecXm+oHumpB+r2ViQBu84rvrHedg
oE1wiurK+jVIaAgcHuRTGwU2ZZv5wLJTjOtQK0Ta2XGa/TIBtOTeoCVnQj+K8wUm
69DiC7Yss5p/o0Ed/kUmbr2nsPCRcHjfYAJxkk53gDy1z/6HBR/Ggj1QyNiPPd82
Iw1tkDEcxIxk7/63tsPDNcIRrqHx0vVum6qOvOGBG/P9Sxy4Ll3PyQhxE+YNtxdP
PJl/L6wNpWgLuDSD0hOk+FLXkZyz0ZVb+BGxhNOgzTs4WfgHjRaSoELYaY1aKMKK
kdS9TRAKgvg9nFZDFsRCnKshf/uOkfazlzdtBlS1E6v3kK2w15K2krTmRUXm5TvX
969nigZhGGkvvmqxFiwZG6B2B79JyEpY3Z5beUpGz2ss4ds3kVthgQ40WgWXVi6I
/i5G4b8VuY0Ndqyy3QJlJPEuO4zXbONfsFnriOe9WVs1Si/213QNKCXEJL/4WAaZ
riCylhiMvxkkdY9UhQUAvxsG98BxJ3Ob85t9FoSSaACFoFs+iiPTql8oxU8hrBJQ
chdn8K0KlfLshbtQKzEjleSBN5PoUJVbb19zDu9qQ/kZBDnCCG2gKCPzJYUySWeF
45MjtPtm9F17/73VHkIpAGklF+MFQA/oRnK2+eZF1tKlJSLqMTZS9dy9axJB+s3K
kz22949HD0OnUJDEoXUTfQJNX2TO1IICi5/nyBQLa5iVG4zrIKNPH8ZzLNmdh/hZ
Ij0510Wxmh+cRDYP9RBCaGH7OJuUk+5MYr+dwBq+4NOvU7YhTICaqL6lQ7Ywtrr7
CyBzFNsry2KONj8hlGz957Bgg3uxvMr5hPz8hkTNZEsK/Onj9L0tonnMMzpXY1wM
8uCO/nI7+hMF3ZF+DjtyOiiq/twiSihCL1Pqn/5kqAPzbwe3fqlkPQS8rY5THmYU
48zYTch+EHoaN55isb8aa2tzDkLaNgR0J5DQpEgiHMtV+txJVkc2Vq4B0v+CibE2
HY5rrTOkm9XAgSkChtxxEu4vaYDfW4ULspGiVa6trcby3Vn+Si247lUO8wE0x7oe
TXXXxq7ldx6AOqf5QYTod2rJPMwKCmoRai8XsTwYxt3lkOlKzUOtiihgxgtp+jOe
HbDnVihIB+mvGo8lO47D22MIihs6t756CV+ws4gdHbgWaKbdacrihBLGLNpI8UTI
9dEUzMUhXnAzgZ5lFtgSOC0ev7YGffk711hwMd8Emqhbt4ySYh+yH2IYUAc0WfYq
mfc4JMsYsmy3/NfOyZL8W6Krs2u1F+ykxtIzER4wAS423IzdFG82HchUvSx0LKmR
srsZbSIRdwsR0VgtAXn9rT4AHyjQXnjm8jWI/oHM2qaE1PZ3sxGLWYF23pt6yVO/
rFQMY7kA47SYgvti/lvrNIqkGDZJ3/ozLlYEysWNBsn98rJbkZZIwE5fpiBuCK/I
wibVGeWbkME8jwTaBAJ7L2Q5ZV8SKfM8ChSFoZ5n95ylmlnuFUnMFsaulTkImpih
i/YIf5+GZMrQuNUfa/n8MhNESyVubHZs1e7hGTedAcIJipx2QscYcrJ3j4xki4zM
Ln1t6b9HiuguSsN7vmuJU46JcpR7nl/lvJ5J+eoeLTt2VGU1kk7YnnT5dWVm3kIR
tR/AljsfoK+kslitjkJuflMUbnFVbydBvQ1GSq1uAUU1zxjiYdIUBeXLaRsOXpbS
splb5acA1LdMgrXRQldNa/ZbwIpvXWq7VouD/y1xvrY/U2IoqquScdok4VPql10v
g502OQfv8p7uPnMM/JL83ebXu+O8u5cEGs3xKHyk0fTKy/mwDxAv3J2t5P8LINJM
k9qt7KZXlbWbHaBdUE/TWjmWN+gddr7IVXKKmkhj/5YYocqHxVzaTusUBrukatXZ
n6hkUMApClAJPF2eWVPjcvKnORD/61QgGOdi+EsncvGhRc10xPly4mQBzc5Xn4a+
UAG0axtnpcGpOamCXu8i7bZy/SZ0lxCsqbNyaPwbsjfmOwFKwmcoFug8LTF4ole3
WED6xuGrWC6d29tbUjr33TgBFrmkUAjFKU5TiR7LOfrOilut5+T+z56CrWd0hz0r
UtGgMOm9BWXnP9EUbzUscI/kizBAkLB0iezJHwJ2dY+hgRn5XXRjsM1SfQrmuuJH
WzKgcCPRCVbrIkFpH4vOB9fBLCMJWFH/3JZkmmxbzp7oCY41ujFd22FOE3fvGWFY
jZ/M2+zbSNuwSn6LjjXzydfwPnsFPluxEWevrNox0b3WIHLp/rJwWYepni9gp0i0
NTcT+TNMkmWmFwMyLN86j+SGAvFHIPi/wEjG/LKQXSATkFp3amN2tMZxkuWrLurV
AWnYT4aIi8EYO5Maxr2FN5Jobpmm1CE/IaD8/cI+Ccwrqtnbb4YxiPQcDNmUT1fk
lyn2PZw6GKQjNHDMfOlFfzTWwS7c8cSyAUjbSslmMj5AIqOlSnBbZCjhnzd2vf+f
lskQGuvTuDC/UZhACOr4p2iTnFLizcwxLSQqF3/Bh1h0yyq/I+pwOHbn33wjPDAJ
xRc0yM4L+ZOaW5a6TESEfxychRCgIq9dnb+PEBEZHocYCaGRcH6DbHltH5xt9oY1
vMl2+2o5uMY98AxsGGitfZhwFGAMHBd3kIv4RRr6IZcoDCHM1pSvRaonp29OYHJR
yvQ8L993ftxU0TW3uDRhXeu1jR1wIDr9AwZUQeuopdJCF8mC38jb6eX1jlKi0H8f
L79YVDrxQyLkGCZT8fYZe/Z/5nXkX1o4fuXyb/1BOAh63uYq1f/ODSXhFRWk8YDZ
eGRf8vl8QYmSfszjLl6OQQK2OSvrYRchhJ5b+VYqwvSTH+OcQeaGkYGhCf5E7zzv
AI+JGIIoUcezdFWljQQ1FGKPhZBXOpMAmxE7NRdgudC8bJ9TJV5bK6x5ezt+wqwK
4eQR2AvHd79D/HMXa8MHb5m6YLqufuGucrfw3PYcgi+jKoFHuIDQ+wxeusVAqSic
bg9t7TMgAyLO3Ue648DgshwnjiFVSNt7w/FEX0zsRfPEOduBqArS2oT1QpNxcBMM
XGawwjo1xWqyxP7ZzgQN9SxxG4vpQjnNGnMXQ1pyDlr5Iybgko2JOjA12zkYLrcQ
m/lby2I39S3GWfVDjWj6PLtG6QMIDF+dQ9pwTQi4qyh/Us2JDbti5Em9iggIIzHD
MHEHgXfvlpJbCbb5/g6ZOrKiRRepcBd67frW/rWvMYKXXu3LVsipu2eLt1aiZPuB
Q4q0Pkwujgn/167azd0HrCOu/x88NN/BWT7M0PE8tMlc0pM1CHB4RHHHi1j/zGTC
WmXiOTk7gdrzqTwBVDvAhbH2CxHV81B3MXjIybV+IOTGX1y+y7IGILhBICXb/OFJ
AhU38Np2MaZdA4SQu+/dCjGVPTfpKde1+nUPL9VH2X41ieBaYR4zamEZkJxeh/vn
SlIN4cH2gwrRxMtpfwJSejeFgu8jlqk5oDfhFFiMi1c3nMRaxmxFGf0QBwUQxdjc
wkiQvo3ljFzQdlUsEXPOD8/XwCfH3l3Q7soesadZidWSbt4t26F/TEgm/4LksOO1
4Agw+txY/3ogFdtTREOZ2D3CYhM1GfpUw/NdktPOBeEzcEV4NIr3wVztTS22KPOX
D9+K7gdPdbJyOg/qktUUVaPStq/TQpU2STpW+xsPRY800z9eKhP1+89pq2MaNHn9
Ebyn5YfUD8UxLQGKavOXSIMGLoKpHVOxonVC0wvcv4CdEm1LXodC4sBGDCtKCKsD
rrne/k2MtSdp8pyWi7issFlGJEIIpGRz74Tm2obiIpSpSjvKC+IaD/PWtGbFj1Tj
uaLNpIbYBUp+MAE9jTVrNxORQLyxiV6ygl4ph9HP8yMiDZG0mL0+Leo66FO4h1G8
MvAJEvtPrT7ojUiVBnf9riYuYovrtxykXacUYePCdo0o/INu5FGNDwoFuYzq7+fI
zMA/1MdQ7kYkZkOmrn9VJbpv6eiJiZ80Ctka2tOUXJSYEJ/uX49ROVxdRBL0xHug
iijswFHRZB9bLqMDBPcCbyozflvGJPgfhYS4m8Fp7qtXsxmQGK3u/vrRVSusxkDw
dVcaoZcu8Tj+7iJgl1Rykk9pCS9+b3OmlxT12ed0FHHxfJoUmgwyUhXj5nx935jU
gP83zlmdcfM189BvqMrbc/iU2CEtBMYNmUZRv2mu7BpfmR4ClnFSkzDopn/Oepnc
WxCXOp7Z9qTELLP94zn2vOo91HZWXLxwgIJK5ZW1VFrMboBOq6SUxIh8hZ8GGThj
IQBVLE+DKR+uuSOxJ0SbRaJpRHRFjZNFriz0THsDxB8QWCJZk0C9aK8Nn2l2tEmZ
1g3LSgGv+czcMWGDiw/qO8kdh7OPUdSP6RR5Xy6XLyipmhB/oRf0v5nl4JDS/rIY
x4GzhHgCiapSXCjs28Vf7A4SwwM6E65Z4ngcYg/s3Pxc93dVPuNDK4oWPSwtUKNG
yuTSkOpWxH3t4yteCQlw90m/AO5M+kb7EDGSvUxM6H/Fz+IVnZvGlI80SGkHUmKq
/yiBNaDtRtAkHjHEkEDjaesJmw8EVWK4KtHoQ3ZT+Gf5GYYTUcGdwR8m8i5nZeVg
jQCZR2eBYWKvLmuXwLe1c33cJ1Lsoa0gZ8+cEYmDjr6ZjpXvH0jIkvojiKmm3/+O
wUcIzZat2u6Tq6ZccrOEXdkHm6U4sMb/AUm1DonYGd+pCc9lYJYiR/g90ryMLrW/
jbtHBCoE2+hT6//wcJCP3LuK0vR4QVTHqENb1VfbtX3eZsDxN5Yz4YgDlz+5Fxzs
Ds6i8eAmP3nPi3pstmk9fLpN54pxesu2Mol5QmQ9CONaYzKBDCo+W3ARqgKubLga
bsmsqJLHb7ZEpeb92o6DUk4RI7oDGKuDMg/K3ixbSmrTuKINrPqmftvHkq+q1rRu
fXzhhu7Y/140kNzret/jJkYoYt74/bCfz0cR4fcU85+1pV7R56q1XpEG2mX7eXpX
uZ7/4G+EWycoyqy9mFT2yF0llcaWu9XeFzfMB7AcAYgDtvh166qAnLz9t74bmw8n
WoTm1PGBOEe+Y36OkrSQykIIXQE/6wMtIffWB/N0C4yZQ2lTOpdCSh84JnBHcpY+
r90MF+2dzNvBR5DBguW8W9ok4mRSxlKUVhuYe49hflK3LfHSY+PsffgI56RaJd2P
N1B9ZaVKaZiMOHghFVq/XuaKkrwk4BfMPfm5ZpXn3SXJqb7/ARquHoZkk551tSJ+
UH93tLK18m9+Bo+Uf7hJVxL6sSwiOHiLqJCA0yn/cy1Li05QI2h1y+rweRdNjU2o
EoUXR4S6do/xhNnxyOjcoI9gj2TDR/6x6XZ65QwnVHmQaWbuRZtn2wgHWltF/EcQ
STW8mFAGkFpJy5XHjsvvhlIuboRdgC6f1o1Vzufjd88aQR25ufz4NLBtW9S4yJ8+
Bil/RddLJrRJOwt/X1VYoKCmOgARyxFjDfhX1ai4AIvvBnp3slW27cJF/+HX4fI2
/um6NhOjN0hCONipcdp4KY/13HnsFkOG5AEr+zylnZ+TKIrg7Vc/h1F0ZeyQxW8B
3Oh8oYUJ4eBDbjm3abQJsHyxk0J/L91rRGURJfA/XTH0rroy/2zFIswIk3x6gPJG
XvUsbzzkQpLxEHeGc/VrBZggmaH/l2ReZTuzi1QkttaW+1YJGLnApghscliEzKoo
xh03Tm/OuCH1tYf/v6E9ERmVPWhdKWDk+gfrOeSpTx68vSHhXQCv0TtcpQrhIhJS
pxMHzBdP3LdDMVP3xaPZZMyqFEZo68eftQa1+LeWaFu/lYVykFkkTD8VH+ckAYCG
0q3SUOcHr6NYQIVpSAfHreXvFBH0QarcPpHvcLpYbi6Jka/akRx1gUc6I8OyktT0
O7+XoA1vWwcNeEYybCgDDDBNlHFiMafGLHr2Hxcoov/lGaBFD3cvtAnAWjQgEQgp
La1Jzl2EG2niXWd6uGUJhqVf6Jri8CqP0x4sohuRTdfO/IeRbbHhSaG86B6C9P8O
UjVydv5+8V9TuTM3DIoghD6GO9vo+MsZkGyugnnMGIuBEc5uXV993qA1+MjXJaxj
qzLRfW8PzC0+oKgaH2SBttRB6phWZ/TtqfyGNBjqy7FrhfBtJg7VWuJUhd0ez4K0
rYZx/RDwDXne3G9ywSwr5lvNuWLOk34KaUSZmhpVVenuelOvg8O83b0B5wlo/UbS
YSL7EM1qASGsq5I0vXeBpvauCSsoGxbq7TREn+VPRRaNznlOP7ChDkueRUtBKDfH
ZEaPofLSmfxcmYAjYJNjCDK0IjIrYpdtLhJgw+5YHQvB7ayMMxc41aodFjsGv2R4
8Cci1n4L9KTCCkpB/XJmcCHEvwVyO1HdA0trg1ehM+kbIvubexXBnzFKYAGdJO2S
vueRegG401vxPZPqk6PORA+XE11/ym+UJ1H5i6m4hwom9mv6A8BFRmQBLRpUma4x
ZLNuN+QjT/9rlSWVHTu/0ydSWHRuXTKc/AY/UiaxWz4dnyPMDuncFjUAhex2yu7N
8qg8pUa5kGVsDdt2MBdJmZEPFStN+TT1IT8m4YlXlvK/L7MQho7f8kbrE6iMSblr
GiGI8rxDMGsQq2yLoMSPpD5ta18QwxXpB9XCK97KAFT9wyn3oe/vY/QbVF0ZDM6p
fE7AjePGxgD8rUQf2AxvZdCo5iH14thh6gvg13Ln8wvn+m9rTXoY7O471XOtcShl
nyWjXkXBMZUMIm5GIYTUXpEtoZf2pisUPJNvfis/1+xUn9SJJilx04PgcYWyWXBN
QSpT55SjPfkYxMxwPzF5/m9XXFc7Rq8OU2vDQ8Y25l+w/rm54SFICbTyiMI59dda
WrAU4uOmAlirVj2cau2Hc8J0m1yw0Ngz9IR0qddr2ysGOOXtArlqQJYtsmn03K9z
Ju5p0qKpSdcE20qCo40dPYTi3ApxElYPMnBT56iN7s6foN54+qe1lc4hOAXe1Lto
6EDDurTVZPDYP03SLtQWvHGiKKg+73yA66dsFPgbmaZ2Zy5ztJ64ZCJ/wN/s06mJ
ETufWb0j/Cf0JyXKF2LsVn+9Gc6OtNZ1CtUeL9IhtlC3v8DSjF3umo/kSSWJgAzO
s7ZH+1/18/cVRMxvTQMUSqofmM2VB3M9MrCpNsdYwzHR5Cv8x5/KH21jbcbhDp4c
PmdUswsRKqESOwLV3CPk9xO0MDN32HaUd2zq6uozNrTQrBndjY2b0okdy8NMd4E/
/SHgktx6SPvvluARBPAv32QSLfleecdDCE+IrzvPrGgxI0eEOH0Owwz4xHT1gbSm
g4Sb5ztzVaKQNGVylD1tFp9VdqDTcSs+X5OEpGCKhUCJwYWCTVwFlEllDs1idkql
hX9pc9K0ZpHl4JmOnW79LsMLjGZcScWz3BjjSEtFqy+vFVP9FYrP069yYAS3R89s
Js1uFcJtsTNFKyhFyxI3+QRSwbLs6fZNjPht+W2KGxaD1w1R5OsY1z87e2NLRimb
eM2w3m8pEQ8wNZQXvZNIk2skE7sgBRfQNbs+Jd49m3sQPMLXsfX/BfQSsKgcFsSJ
1GhKbe2lPiezljSp6qu0STBFZztXnHqfmC8f1aNm5MbktuV/9FavlKSTGKkUmMwo
kf9MrH1pSDS6xYN04FfeLuMB3YweVrKEwU/UuB4uriCXYIIOSlFEU58G8+6dUitF
LFgi0vlQl1s0kGkCb9G6VGwhf+EGJ6kmqdPRyVuEnexIM1arR0UjUj6ytVllCEIf
MjJ/9RAHcAm2fblJxcKn4hnCVD53BNaTKxH0gPk8Bxazybyrzy0FJFgBFcN1Vkzs
AzSZILZjdR4YbMyAzv+l3ZtoRDzpy6WWv/Hq7Tw8AttPKF6wfslBmip9QGC8aBNs
5HM645B1D6PT3/mSL4Hwhf64bKIx1VYLrYegAvgSdw1X333Ac+Mn3riW/Irnd2ST
DA6OMOtWxRqw14iUfgJul3oGLBiorpgR/hwNxU65FTjiycP3TJwQ/PPVfmjvZ1Zu
byMkwGBV0Kz3q0M7kTBMyXH0KkuIvrt9W7I0dbmgbbNNl3NZk/Mfhm5gb47frmch
PMPKTTRoXdnfhUsCGR1HNFYFQy8sbcCMPBBKWmrFVrmSlo6O6WfMXcmgIGfe9YUB
opLQVWVd/VyhRcQHOQlAvQwmqLg180KzAL6tC0TlqO4QKEeZ9hM/F7Gx06angqcT
Gts1ODmBnfxjk71+De1NJ56ae8YVQPgK0Uig2+RXFfyY4BzJ7nI6t7pzZDspgYKH
aFW+87QiFTVI62XCHtxpqBdbcbwdPDlEQAVrrzzhpEia07VBZf62RJ1SykT2InjP
zEAs64rp9h3Raz/dpWOLzopNxN9keBVAhX+aM6yvebjJ6OGCqEtX0ofmCjzltJok
lh5Iz6Bi0YQRVTdRQGUnGq8Oh8z54CJVIwzEP3diIVUernS1kAdkhfuys+UJAPwG
V8tGWrJ4+1yvcMNzyhkHXVEoFhcLJLjWvXYa/mrxAHA92/v4VIQW8LoF7WaXL3at
TbQggUPXY9BvqQyO0+dATwrStoTD83KKsyO0sJOY/M7gIXLYooT1Poz4S64KieF1
NtTr4rFwLMLvPnbPTr99kBbTM7bIXgPad4sEPieHgz9xd8Qvr50Ng+E240onYhoS
1e2vwNPMv/Z2LBOUKpp3i9cRSm3EYfn78yzkeG7vrh2ER50IUdflym3ES4vStc4R
k1TfCu8VVB2raenireZ2J/bx/RXAw0SUGOCxTFhvQr9XPu5TST37DMZ+Srn8cF+v
tUm3HKB2dXj4SC3euanMfq/MESlpEwgwumvvjg2u7BsSdyiXuN0kxnOTW9h1c7ya
JQlMccKDYa+OWeNlneCZOh6XgtunPiMN6Ml7c3ea9huR92KFoRMha2PL3x2cAHMD
gKZDXAe2EoakdcF6Hsrr0voReqk/j+E0ZnV1gis+SbvWXwzrfv4mZHbfXkQG8FDc
YdMe4fjHNMV83yiBRyl/mc4GNXp1tk7yXdNk+TmIzh08YJwLLXyJTo+aBR4F+/s2
HlfEq5pBxhFWuylM5J52bMzQMdH5UGXAbcT4lGOf11+I7h2cL7bHBx7cqQAixrJr
KiOWYJAKn3kB4/J5LVrvtzoxVUiUhrBgQCwr1VT2UYSfTKJbKNLI2UBw1JHpfQls
8hu2v4WtWHribtJZD9MVuzdDN9YsVl6ephtNXWLzzQpRnkF71Btg+FGiX0ouErU9
OzFDm7MdUIjWhUdKInDmExRq019p/PEvIgXRgia2RLF/ipGNnSr50uNCk8tohykX
XcuB/YbQPmGU+eBDFY50jfjTF6CCx9bMVmgAyFtCGVDWyw/F26enXRFqlz681MMp
O90pp02ZpDpoj0eOj8Cl6D4byQVQFDKZ8bmGT2kg16gEgREKBsDxUc2NTL50rue7
l/hVByj2eZr34hrHoO9x9hldh/4I2vjvWQEhew0qpb3L6rZM26dC5IwIiiajOZ2+
CP74SvL7CDbi663A+YnVgK5JSIhPeeFKpXnbzBttMLXVeykkvYxz1Vo6ifzJVaZZ
6L4B9kEHAGCBQoYR5jQYySBzioY7E4W1aVNuNQDjZ0XHqY+U2bNacCVp8sOupstb
Y4Px9EbWLnGC5BQeaSfNECUmdqcoC8BitbDpwBUM/Jdn8LA8q1kX93z30bEJHFSj
24lXEJxDpCb1lGCEkENjO7zQ2CV89dTfgWu5/1DaOweZ7opxp4OymDA/VJ4KtQDc
dZPbbLnb9rHeS4UlmJD6TnBsodcEPW5FeKLoaIhT3kAd6UbBPMnm4KapxfOHe0ni
3PNF5KCAPwJ4bhp2lUJng8fN+qtQgFlqUvNkYOiWZVv11KPHM7tYzQfNApROL6hJ
F6ioE4SYrc/cQIiyaOxB/EwGV6kvBNo3Jpewsq+ivx1ksbMCG/y+BIRpxROd1QF4
2ZXye76eeihyE+vy4dqoFD0KYGMwYDFMuERjSEU42QO/h+/D1JfTo4U1DUNcbra2
4NN/3talIkxtLkv+x1it/OaPqPyX84bF6r2Ev9HdFM/miNANh97vAlvJ6gvYVku6
3/qUDtnIjCHamiIEUz/Aj6RAP1Gl0H76WnyMiPWuo3VlpZ+60VTWs7dDuMrBl8Y2
wDEUpMLRVskO6xY6y0wpewtN1e1bwfu+4nQzRp0G8hfrTyVgpdwaoqyV9tbcbpaB
op4o9KkSINnjb4AmCK2YpEceBV7V7TSy7JVS8k+oqgHOiqK3ulQMqbyhR9x337zN
AcGNT6QT1cGUAxuknA49JZubs5bWwVZpbJmdiJYJ+jUSKgQBOXn2iyzYA4q5GJ3b
yCrCED49UQBcmaC6+3ma3stY/eDOs7CL8h8HuIZa1sbUsHBIxmLLf970gVVy+FnJ
HLIaPHu74VIpFls04LtnPaMlmgYzC3k8hGy+TR2zkNr+tEadWM7vtx3JC7OiuEyw
40MqZvW7SETNLShxh7dkoEonr1zdIW/33VnZN/4+/DOeb43BlgmfyxNbCC71EzmK
bFOyMpvVjEycbnnXtnO3Tk5gm14F/PYK8XIngQ2mndbHjyRxED5YsGySnc5p1DWn
pJ00M808kWZSTDOpb7bpYQYbfcVPnZi/Z36TcX7VGTKaPouRQgAqQL1ATInM3DLZ
yXvtSog45ItotbV92rugu2IZ67h2FqdvWG8slxoMqt+v1Hvwf4NoOZVtIwpIKbDm
1PxFUJDX5ONDUVziCqlPR7K0LeEZdDnN52PVqNPZqyJbtb6e5orSo1NA68RD0xXO
zoSiFpMI4JlRyRDfdgtlmc9hmBVdjfakqBPR8sgwzAKoEb1BYLFkUh/FMLZ9kouw
AXSDg2T5FMN8EnnrJFbty53ar/d/Pv0Kdoa+V1NEkhQO2OXNDQa53q4u+QCcLTcY
spZG+iVoWaMdMNfpQZ2AWGxPcMs+zCx+NR8Jxkw1HDpfBqEMv5I0cNfhz+YPUiCz
4/I8GprAN/jW1i7TOdpe+/qI7DS2n/gH3OeY2fOhC74GKwUF62iN8nxzYQF4wdQc
Jq1e3ki1/HGNcprNJheqmFRWInnGtCmMQqPxJJWI2y/526OvRcZdeE2ha/A9/lFu
1zRLbu8/+IdhzN4NzjfHSIr3NNRkR0YboaFZtHYgCGzUPhJpin3J8MNo+lScODnj
P4iBsLpIel+BvpS4K0kZvZrybMORzqx1E+3AZ0zBXCAtosYFMgqrB0W0+Y1xk/Nk
KNnXtDaQ1r3LWbk3sc/OYvSB7wXF32MGznGwpd8mRDKmT9buXvFqo4YwxdlNIB3D
hIbLanLGDxo1Z3OhhR7mRvV8Wi09hyPcgy99crw2E0uc1qfJiXdaOfyfm+f8Tc7s
txFLAFYluK0MDHeIV8u7ZxDx4q93vVNsIa/Ra0ZNYOHedVGU31d5u/Kq89cTQhhD
/FwxNMb3OuX08pKNyLifsaJdvcwLdx4H50Cn5//WG2BVj3ajNCryVzFr+YK86BHg
q7JHY/g6riGyPd+/Gkcb3tUK7HHeXkE6FKhaWgJWKJD2glYCf94eKiepwItOYOwF
vz2gNs5VntVe09YJZQEnBTpElGGZx9U3SII/UqNSrY7Dd7Cw655f1YfP5V2dgHHz
uPVZq57EmHj593Eyaj/ntn+ZYnSos7SF0wfOLJV7TZpiIV6Krmt60p/6m5xTyP1E
qDUN9TzE8bpls3vOFgOstJRvE5xndhUF+cjVstemn5l0LDCLhq2a9qXi/LgPiaOC
OUOF190rNno+Bwes8CG4vfpjVgHvXh2rhEFqwU2nDfZyPnp5b8kKOBS74VVj1qVP
TEC4mPvd+87jOWg3PyT8dcyiTjHLAOsBq0CzJiDP9A3r8UbsQRUaFdH3mAhPTP/5
kYscFyLITqIZamuPgaNKUhz8DBfrwRtFdp99Tuhk30k0TTyxroWJHSxYOUKPOuh3
bN+wh6wBDA0uO+sQAq7zBt9669GCVf6ax05ThKuJGAfSYE2ck2IMZCf11gHCgNON
AU+hx0SFSamicCeFO5bEsbIhSFXknpKbVEF+2e3sRJy5V8Kqo4ezUuB7dJV5sBXG
hkE3az2lG+GZq8UfzreA0R6iiIeQHbQq+rcfYApIQKUyVouTA4w+JJLcAkA62q8f
gSsNR4rigBljyHrnED7rTbg2zO15KH7Jcfo3Al90lJVlvRpI2r6c3YY/okuNejoC
RoFcUHjqSx7YwN1H4YhLTm64Mfr+go5QxzQ5LLdLENryqEFN0uFhzc9roMWOk5Ub
RfmJuNihrWz2UfxPRHn7ZFYoys217IPqluXgS+/x07tlUlBHo/X+NuohrhceKZ9e
xMUBk/HmI6iLfcc5MlOeFut4iOxneGnX2KW2Yj5jxw3BtizUHNVAiLdDh/D7anid
UALFjN5gIet0rdz6VvfAHCLiQOOx1jEx7JWeJh5hCjIIwi9DqUiHLyrQdnBTc8TQ
AOrnKolETnKSvyxGYQaNHNYr1SqXpIXrMFeoEvDM0+n4bQ59IYWE3mSH49p/rpjX
5F/79yFCYwyOwTEOuBYvEISRgaKr12QApPimyt7o4Ze9Zynx8jlUe1uzNZtVPQOB
Ae1bPbWyOik2ddlVOWMbx985MHuxV4RYoP29ZKhXB+qE2YqYNZXHGtb84dk96+WN
GvalnmIoGlYoIffA6LsaJslV6sl7MkA2kUCkdNjA6d+GIOgLMg0kWvtP4q+F/BVE
jYC4yGr/mwk6XLmxbQ7h3U66GZdO1p+U2tvDhyBLQDzSmJusZ9NJ5701QQTMs7JS
3nWa6d2mglv3tpbPfWjKyBZX/9gZBalP6vXhZ1p4c52fTetltZ2rf9t+g6EzvwqB
5ns+SIdgqK1B4TiVwfv7c+Q7FKZuOzUUTvcn15LKD7JMkr2c0xmmpUrFqRO+UstT
24/ygOuSxL/EtIaaDo8R8s3muBv22lIn6sq9ZHMj/pnB85OcQfA1V0m5iZtb9sWN
r6d3fsOzpyTvZqX+aGBCDEi8GgJFucOVbmX4wB/yk3GRu3PxC+SiEnwwz1pk9lif
lBNVfv2NKWJnz6h+2bLEcyshYYUJGlU8RwIFZ4tc5ZGx6erLnbFUCWQ8MhhMs775
Xme9c/C/lMDZIdo1bZjKKZywMSJgj4aAIDcZilf8UpcAzDZbjYHp67MLxaGX2kJA
0mgdNgcAG+TNU31cduVwUa2cgn6Swpg2cCWo5894Mi1DCMfw1RCNHyKfrG64Epc8
hfJYVp4YwemgcP8+NA3OS0UJvNTnx3GjjZqAzkMB+3Aw1rnd8CL21pMwemJXqyA4
T1uJ96ZFRQrDtr7/MZ+O1KDY79JCxdBqoi5Nv66cP4j0svpHoiPgsNUDI5PHG64Y
Hzl3K2/uTmR57mzfaqgXmLRNsMyyOGDQifLXOTd1RdekNdT7OyBfIG6zyWgKR8on
nG4+yivjPteqAuVOQ7ExfIdfbS9zi5dy810TkmWvH28QPuWIoXhiTzZHpv0OUUgQ
8sQLoSwWtDlfYTF9oKUynKj3Awrlgx10108wopwJgaEKJoQJQIRLIJm6px7VOuOb
RfoGXIDTNJ0yxTG83sZ+H1VTLJa6NYekGq2vfgTQ1wHbdv353BLTFVjwS2fD3p9R
39FO6J5SukYz68yqxdT8MN5ZMwW+Yz1db0FTZfOS9v6oehacJ6H68pGORzHsmv0B
JVvnjxqCfpyFVhIz8j7FXW09V1f7VLEnTHoOSn8U7XsSSc4hyjz2zV+i2e9Qwtrz
WXclV+gGMDGinhkCiccAAVdP48Ox2pGovK3qSNzWJ5obnqr4jwi9XX4l8DfSDs7e
Q0MoLwynuQaZlHA/jxJmiEVTApMaOsADedoHOjvNwtVXFmgD6X9Uci3elG0aKiBI
eCgSCVIqvq6zCvVjhZTjR85AMUYqk2hvi6vmysU7eq+zIT3bUMTnNd7NGh9Xu/MT
grNCI44lBdjD5AZtLVUuO1sXQYBilRHAaGaw5dhp2tFVPhAQ2iQlpbki13t19Apg
mFwP0rckrjX3caqjRmbwqWswl+X9xLVqCNsED5CpAMWmfo+w1tb47+ZIoeJo8Ff3
kZBQx2LpOCTwpIirv/OwAikV2KKr6E0EAGY8SxIMQDRobC6FaZN9ZxvoT4jgW7Ye
KtlV92nwCC71ZDoDiRHMBlDjaUuST8W4ntiXLK3Xk2U53zCqXP9uFrHG2dSlhDne
CPsI6Dkg1mk+eMfue41Ri05t47Z9v85d0xIDBh2yngOu0ubnnz4l8UOcGyRV8t5x
UXGSjUGW/qhE8Ov530MaveLKzbSHiBRELLdKEbJJG+0T4HhWswz45nFEci2y+hnJ
37WxI120NSZ3M/kujZHpl0L6Tt/ogA2MJILLK17T4ANpiJsu6w+hmQW4oCrOWnUj
bZz+2vpAVxwJTJmQQylQTJyYJpq8L9eHlgAak6Ss6DoYtpPN5cJYlYKUcvLv8axy
Rnc0PP+JV9fnBuknM4i0gN6BP0xON0cfUxNYGWPWoGSl2Ned78m6vA1zKCPLxiig
mmB8AScWhbuw7OZoPZnP8isTlQUnEQdUnJ6uD/5UqNsDTvxV1xzz87We6miQdp8+
A+CSJJ/86QkIOJRvZ8kdgI1VfHx6Jz2RQWOxBE2pBRmIQLRe1UBvUlRTyeI6DGxQ
EJTRoWeYdhOREWtVAI9rbFSRWUNHdU8k5ndoKNKcbi7FfbPBGB7vgbLKG7FDNhDs
D+IdiLTmy/udI0xs3gGMfDOStLhkfjZsDUxMGWHILwsZBt6vRKozR0L5OCXURuWa
5YdvZNe4Yhtb7p7BK/jKuV0EeEeGSJkh2MvlZIBZoaxc8iNGc+jKwBaCjpv/0txU
FAIJk5ZRgSrfq2UUIsXIoUrDNHrRlvk+IVPAVW9V22zoCXw8xqEQ/TubY8bBgN7P
Fzyrf355ke0FVmMSSQ1jnfVmgRafRFpQXFUmBibpY71jrTawX99Iq0jqRtsPFQga
dJiv+THXDE2/6VctsAHXew/8yJ05IC5gaFEkXw3pI9t+CqfBA4JQaGxI7XRHsJxQ
NAGYnhcoMwaQopHI02inbFKP3+Yczmk1kYjZghH8gZWDATStDEyegZwxMxtjqGLE
I8DgDGhkZ0xdl9jYSglHAdf+9wl8m3q0s6jG82OlIqm0w//7KYHZCpxiodRXNIWz
frO05Qhbidc4fgThMnEKtDmER2B/jrceqeuZtt3dFXWOzrcCPRtv1N9AlPnl/1Pl
AKzlvmdpVm3N6hUm/ndXsP1bNwU0XY/XHx8F+80FvIckhDcVGI+LkuIQ++dJzyqN
MBTe4kBolY8oylDcoDBBLHYeJrZoiePJKQyXX1rD3s6sUG2zGahMi5VC0HCYbwb2
gNR4atlAGeY/ih4Nf9naxX5Uc1aW4vYOqTGR61WeTq/phVJJ8MLckQYxvZP4ISO0
aAtM/JUgphOio/p0iOV86KKrHgj48q94qsaycTorXaL5ZD6Iu/oeCOz9A4FK+SLi
RxMjCtycZlsNcn2FD2PDAQtAN+gOR65GjPhduOD6sYwBiLrmUpQ3juniYO9NWh8t
BUpDdG0ium0iuAeUpnxCb8DDV5uDyPsgg2/7lF4a16ZTkO98mvH2k28QQi5bpL1R
qjhwP97+NsO+NkarzXtPBpYmoBtem6LB12CFayXGSESrNRoxkeKPS99iszR648yP
nez5tqbLtP6C4+wZNksKAjbxb04qdH3+z5VWAHl7j/aVhrwTD8uhMXtTmXwQCUkm
YZapjt0tUmGvfKRimWbp6wLcyUSXpTANbFy9dyIhN2NVS4vKNv0GzKMl8e/re+sL
YiSEr3NC8AZwQuIKt6M64VbR5pBhYdpbbjCM3FJJK6r+GwHJPzUutbrp42ojute2
iAKDDZ8dQ0KKicmrbNri5OQJnpRW//gOA+hgmku9nwxjp8yOD32wDe1uWx5g8dMN
IveENYe1J87mJHNwPXw6+WEwvpWVxb+JytJbvKlxbRCAzP7vA5ouUlMgRC1Bu2qj
FqcFVUw5O2WMbucMiQ1+wRb5Z4FTtDQAxfKrs/0Zrf9qp/P4zIpYVQSdgwFRl8za
oPyy/Hya3ZOCIvVni4h6ePouw7iLMNt0We+ZMrW6OlVIZUPrrbQTxXF9v/gIle+o
it1PXZ1IUZ3wjQFygmbiDuz0psSNaaOBAVtU02KY31vCGMouNxI4Sb0r4kq+Ch3K
EeumwmHCn4IBPcZEDpdSBlVOWsbFawQKEGNH7JN2BrnmVdSTj1hSq1YfhNxAK7/Y
7yv2SWv8JxVLlz6h4Jl5RnaEKDOmab0/tp/tXs2Y3Z+lFVrZC3t3gpG97oNUNc3M
EwII0/P+qBlc6t6z+7+e+r2Gwum/s9D/w5IFIlnE9jW4uVJqt5sHLPWfW267Vnxm
Hq10MD5mvVp9qKq/GegkoVZsX2zaGhh9iu3Ia8U1qrLvoPffODJkhnKbonzsy2hn
9rBtDutcYPb+Mm+CPzFu4Q6GRI3faM7xrQX2nrr04TOEAn6H1WUeAfmV2hulP6Ob
Z6BezbUjlN17c9F2NkaIg044Cy4941Vt1JtlVN8ASA+suJpv7oMdD9PBic3g5owk
+rZQCD3V8+q+YER3IZV28C8PE9Cn2o8A+4Khk/kG0UH4T7ic2NZsPsz7AX16ZNec
uABc4EdcMEEA+BEl6s8KMVhkG9QDziY28Q4k4Wldl4kNcqPPQxJbHvienN+0gaMS
AQPdXxYELHBdpIgghl5dbNELoJhUOBkadSC/kPjoMOwLG2ouKVkk06yXfW0pXGYy
1uGAHmYLQt9MziRUd4cGVnlyl/G9yk1p6w5MztS65UwGyWB3iclr2xwpce7iYLGP
LFMno+OgoRIGrPoWD5SKq3svhRQGVhefh0oV5wTlHZ1+V25Pezg+vwNu8q0ejF3C
sxFmvhFE+HYayPfn732CHaSE89aE2OMthCzeJfBoVTjK8iQh/Uvm4h3zHns/UOlL
nltJ87jNYUOnho+1Xzb72xSZJ8LQKoZfPtEK1lAvJJi78Odcwb33C2LT5iyCwS/4
QO/Ny3AsTWds6OfruzTyfPiud/pYNIQlrHEOYvfvl+jLw+X41sPDfF69xHoJ0EOA
Mxi2DzmUAk5CV3yt22aCwxFU983R5WnC9+mFYFIdAvyBoKi6irVLMouWQs/7hQjc
X+fRpaHg2Ef0TLrFYboLNHaXVi9mzKH5YJ969hkfq0WRpBoRCmU0Ez9yC2DFUQK/
JbgWK8W3juR+0jNuOzMEehLZuYXKaplf302isE7ooo011j1Jp6xpo/aFt1zMn1D9
/JvcSXkYcE1GMB3h/bACmqamlGxixZ589ndZ++8+51SyLShkOGAJD4EDBZVNkhZ3
GGfRCbkUG0+c5DP52QkT32ae/gRLRCg3ZF23yuqY3O+MgNjIQCFM+gN0zk/Ru4gx
1N/VMFo51roNx65tppA4J84Waqcy5P1LVvejUpMASgAwevCT2k8Ucq3rOgC5BsgJ
EXSeMJ4uN1xE6u1t+5BFUrAAkQ8NYo3Aooh7oc4C5TITdAEboYOyl+HJCSKbaHhe
jO/8IY1mlfj9VJHRyr2Z3OSM8o4MsK2nJ/mgvMxNtMd4v+SUd6YCsw1MvE88ZJZe
/v4TOK/x2ui3yPpmXsJdnaVJshUtp9OM+QwFzNKmNSNipBqdTd1h7TPFJ7g7lz1E
tgyiSCF4vEx9TRzVe/h9rPQJ3vDfdiASmYF6eSAToOJILRKXgaMwKNPIi6gnJl4J
H0oYB/qXSrsVmNba9GFvfeqN9XciHEQAahlFLI/470bwTp72zYVkTbt0AK8Qpac4
upILw3qbXE8jekDdyHXZEqSEshRxjhtDQ5pu2M2ZzbpHhuvZ2LQ38yMFkxZkSiVJ
dyixhcQPP45bQ83vyXZRYjEEFqp1X26HJpg1RWYiOlOG+K25zdocdRvLB4cZFgNF
ENoC1l1fCJ8sWM70pQJjxnuyTGqqy5b++vZZSuMM0AKVbPq+1SOHDlJtC+8TPFbS
JZRwjJDZLk/w9AC1yepgGwlPr8q8mHuvHxtrI53ROtr3CCFdBArezkgTlqOLCpcZ
3WfvEdaQt8vQOKHfgTRbThP0Lk3ep1NyjW0Tz3jt+Zezr1ejEnjgfBCT2dZvm3jN
7D91zKS9vL2QVlAR6E/37hXYb/E4TtfED1IRJc57Uu9MGey4J7klCImuJVdUoXP9
yJv4GbE/2W9tpaTIFJ3xbpAoT3pegOc1I2HPSvLWLcs23cw/Grqsaf3/haZG93St
zSUJn99cvjROJhq2mzBR1lNSXK3K5J9ZaZUnY2pMXc5OuktfP9PDsFgRcnFZ9gG2
aY4rAo5TvrLjMO4IQO4yoFpPRFc7+WZeClE1BMgdHDyro89NytWR/f/DFHyf+iqn
BUWAGKNIENVvVjaDjxnwt+w9l47PmU5kDuz3dECFFX9y65C9bjB/Ehs/tFNp8wmh
SuhO1torrh1e1jwVzc7WrXKrByOdRFK4wUqEU5Or5TyVUP3tgc9JxfKQfrVJQ7E8
nNXHpi8kbWMk17Xbr32eR6spKlPjFC52wXcp3Qfb4fnzUltqcmAh/XAo4EpP2dpy
NMe23AX8iNE4v7bocJIsLlkZPJz516PBzsDld+OdFJMuyyP17L2irXI0RQm7qL0Q
keMw1GIlYNfCCZLHg+Td4/wmMK08BJQfukHDw037KLl3i1RUjSi+heAm1b1ecyKD
Lhelu+qX0Hbd+gXBByTN6K1XMlZ0a/FOiz8HYfx6GI8FSxxBC/1E7XtrVf8yfBTw
7CTQs4k51KalxiWoMT9O1/IwUIHu7mBllji3caZi0UeRmyne74UrNWB5EhH8Y7uS
56LUZ52mXbWSS9bHSCtb5oJsIe45Z3w82br7TlTVYMBnXShNMnIQzXWV2y2a05Im
YlNZk+PpMMchkLBJl/bwfowfBu9Xir1a0rEoXqpzxRibay8SbDP2tuYZcSehp+PZ
p8X3Lh1XaFPH7nma7LdnM+3gX1ea2cGUgPZrjHJIA3TfXci5QarotqoudA3+sJ/4
SzW9Z+h7F6R9HEU1y4tYiIrvaQ5zZ1b07SxIgf5tuevkyllDmopRkBf0TxChunNL
WCkTeQ5PD026gU/GzqQfTPWpqE1LkwaJRjWoLy/Y9VCAm58uuh2Gigvu9FgkKMXY
0s1h9E/CPXcxGERLUmaiGZ+N+Q3GVHGfLBDF68YXoJWMSeGUElj9BKUu75t/mdOj
T3FS5eY3h6RcFIUJ/T37S4BewAK65juoSTJYqEGyH4B1pdnREks0OV6E5H9wGehq
hkbj/YbyQlomhxPcCJW0tihvTw6hvCXcwAMh0epl95kQNM1hcva+Th2avyzJxcO6
6MLjE8eyLDK5eUwBysljy/Sb3vgrfPo9mRaWmAVizVi/7e0GZsZJZ5LvaFUEj2U7
XwqJOddQYzgj5kM84AwVesavwXkQ0bDACJfiFGtnGH1zrYlnP9sCuvj2PhZ/XT8F
R0zoWsyLB1x1ECttjZZ/ZTCKgX3EA1E3F2SRmmmpm3iulVjsh1VqJOP+LQO8QXHz
D7hEk820wsGEDyevmch3KZsK8tLwpokjdQg5nuycSWGRI999vpqjlPOxcGrtHAHO
aRAmLi4oI0xSlmo+kpKhqkZeYgKS43jrYy0dn+BoJ266QOb91rRYOGNfhZi9WDCp
TiF4+i2X0bPMlzvjRNFsIr+9s4NVK0hdnJLD+88K2hZ7GodqzJTbXf5DILL14G4h
R9s1SOHzLjX+kSbEX02g3L0EqnOz/DGT3J01m66CUVtoYp3EjJ0aR7aZvFFRuZ/9
5g/BJB+BGWB56/9bzbpWZkaCjrUu0Gje3w2QLiZuMExdIQUxaz/VZDqoH5Xe3FZc
aSR3V+ToSFpZBJSlx11/cJCufUsr9oRLkQoMUao3VgaE8r6IgAmtsYz+/p67YWgV
rlw0nzfu/LXMmSCNlTxpi29W2+H5rzguKh1z/SCM/TSF6msLJVkj1Xf1qV8eYbDJ
S6vl5XC16BFZR9IV1zcyaQweKaV5atKrpFlrIluU5OuYMLw5FOmhMTl5jtJmJnrk
0RC11+qbkQLKDr50QEVgXRBXHpDm/YRGcTBtkYDkfoqW8Xu6GBs1aJPlojYXoJH5
hf5mZLKzL8Le3W+kUyPXZWFtRcAGgKYiszhHyv/DPrSyjBLd5C+YScI0fGcB5ViC
GFFQEcWfdvUrDVnIjlvgM8Z5PDxh7e59V3IALMnxNcSshp5bIAwQiogNuPrQm2n5
LijYXq3/Yc57BE/5D/YzJqoDxPZdE34ToFMv3pC68Kry/q9J/XaaAirpKVjPqLop
TyQzi22LcPvNkGiQAhaFozro5tZCbgvKmT/sxAm+8l2s2wA88ZihcSjyyeYOtYwj
eBhGdFk2uwvMGEeZXC3YWOKvNip7hlI51lW/NEOZyxS7j3aHijn4Zds4Fa2Sn14W
MF6j4z6VrrZipQC53qykdQethjDcHOA7eM2PlrgoxtaYgPYtuq82e+Xa8I+fHoK+
xfU6i6YTLhlOc+EAYcN9uvSDqAMRGC5UlIFxVkxX2TchmjtzgvTiY2cvOiF3DZB0
ePk2PQzFZoA7YuJsnxK4MaIuwDyhqjrH1qWtBKGf/czznPIkEFa64xKYY/vyHk+O
8vKUy/PWb2fHQmeYa7G/iChwt73EDnyjwnQ9ZyRvoF2S1OXT4BmB7DzQwVxPFXVD
B6/zbQ8KWZgcki4T5qm9ISggZuWnYfo4mhoLiQOI6NtJ40ylaw43s8ed2sZvXg8m
AOAmvafNs8Bh6bGhS6dHF6iHujRqxnbnI9Jm2kVZniJi0Unibd71tXk53s+zqx9d
dk1ilOFG5awPw5Ntc8/dkUwDAO0pzh3CNCYoUkSaYDJ2o5z3AnLBkOI7rsEZ/mjC
1badyIQwURCDEDaWGrb+2c+sBZ51sYCn+UkZ6kavr9SVdeHc8Demt7vM6exdgAOU
n8+kPoeWDOBuO/CVCYILJSjFGACMNm/lf03HEch+q1uOffdGGW2r0tS2oLEl1bbE
h7nNMmFxOmnD0hprO4VvMYEGFN7uBWxaWHW34vieeJfBH/WnleyYh98ADefONEy0
HzQJsubotsnNkFN7U1ijUMeMTkag4Zr4kXpuWjT2fEp1IDOQf5CPzw4AO+KcLn2L
T86UEi4SmhLUobG9c+l5fcIGFxhTt+/IwdhHyekb1OGhoj0+tB+o6RrEN/2L7yCI
mYuB9Gg4YpWgrUz/E8tpe7BSnI2FvTreMe8TkqbSxk9uOd4COh+hdawdbW97esjl
45ZgRzOFKrapWqxB2tdb+pKg8VUdlntMGFilYN2Wa1WEeh35xn39+kO5x8cyqqAG
e2Pob2c6y+TeqbhDivy3ckVY1adesIeUMxqJKRRMZDXY+XSk+r7GML1Z92Sp27rW
PM4FwpWHl9YzfuVmMdm5vAziyMaVL04HIGLMTVf7jh8kSsM1+geK99F+pLs8Yew4
ifNGTHqiXzbDwfA0Ab0RmJNgV3fvGV5LFyNssGf9FLbKSbMAVXohaxYUIFu9Yy/u
o3sLx4VMQd5lvya35hUeeQ5uE3wrOiCelSBIWI+Z33lFg6DC2eZoMOMo74IeqFuE
v1Jvzx7+apYgmj3zcBQXRiY02HV8u7UJwLnH02SGwJJZP1nr4bCq6yab9TaYJMwl
3Rz4uoEnhz0/5vy1rskCfgH9Xpy1b+3OEuKwP35QV9BiH1wgBN+J48abRYAz219h
OHYXynf9MhhchxrdyMpJvwB6sAMsURDOPL5qurTuZcjVES838R56hjJmt07xrDsr
WzlCeg8P4Ceu4JkBWr2cBojN0cJ+c1cPKeNV9OoNXTK26FT+5FRrzwmUC7LFkBsP
RKlOaRgoE3UmK1RftKWRFWmKxPBTrtrr5MQz1Qd0lzIFc0L95wR5mfZ610ZJ5zLe
LPCVymvUIZYzRB6+kpv4QNz+F2CTR2d2AZe5zRX344/8wp4FpsXNjAY+0l8eNtda
p8gB5Stkg1HOpIaosGOIu9zTTSlZiRezyq2gDsJQfOjv8ZYv6tV7oKxvsX1NJM4h
tkP/AWxIpcaZoYKiZDq+pOjZ7NDBTXgCMbELnl7a13RgVj1XTyozkiPFk0SDYs1q
ysotSuDRWoxUP9a1VvgNXgGYIZjoQlXBahoPRTJl4hNmZHswCRLsoijhQpdjET9X
KNyqJgFDibwZ3g41G7ehn7UK8B2iAUglJMVCHdXQBWNwSiB6CyR/buC13QC392so
qXsxnn88zDr0hAePliknxLpxKfcov496vBiLJkQKqIk5SQMH/VIMMqmFY9VFVswT
D7L0F0yyhEiPwvEEda1n97btmIWLAUxALDS9PD+6J7YP2JT8MdIchiEVGkkz23fb
wHqX8pu/7gt6ONMQGJB117QanagbFJOEF6Z+mCOfTRD3SvtLXVSf8F+v6RGKQ39G
Qn0XNGObvyNpS82ac7GdQj+jVJIriW9AJQkciTMOhb1CzoXYBm9Iv7TFwCgrt89u
JOR9UgFcJYHox5VDaneSa9xjOUos/usIHNhEBc3cA3Buq8d2rczV1kq5qolKlBv1
Vgobk5GK25g6Okr1XypL+EAtSSNvIaO+kGZc5BfYjq54QHxvqB0oZxVPFCRe41lW
5oCgfLg/6v8bLckQejE8aGg9H1P9p2PSiomYlN/BUy+uFmuR3hf4thS2AIIauQKo
UU2JIcLZVLEtSE2NG8jpUUqGdARTGsu0WfG6E6fUSRloD8fPlLPIOkiHmLavOhp+
3F5VCLpazETViJPXHo4EPHZLp2FTR9LuefXDtMIHz6kTnHkiZ+2VoUbQT2KplLbN
UbjWqMbpE9/X1fHS2cGBD49ppBQWxzAi1wu+f3w2Ae919FQzx31ByrRSZr/5sM2G
r9cm/S+xMVnHzlna+Em7Tw08/KAVSFzN4//ZG4i4JKFEIcbtpIAnjKfQq0o7e8/A
nRapdg2MBHWy6UAIvwLcVwqQm3ZjzU7TU46FXOqJ0gHHsYb1KiZczlBUpeFi3HlA
VmLh47WsrER9NRXnk23k1umog7ptjMqdRLc76Dd3CNQRuV7QtGiomyNPb8K7WmPd
b3r4FXaDCxii2d8B2lSU8HFF3yR+dt0tfZaTobhDd4/CSv34vqVYyTCQftbf4plj
8OolX3PEpWlC/tHSjXQtmLML5uGgFXqWH1dH/G+hnwCBk4b4hi9uGLji8cjqa4yT
GnF/ZcaS70IeAK2HOvWe2eZBZUiOGaaDtgmpi2XudYIWc/Rn/WQHW9L8Xnxsga1V
APb3g7Yza7tOKBreOd/TwqHi21jKv28QsOe7cQnizkd9uSPcdFedaRupS/JEx2ta
uewowjcSS7E/5t9MfwHDFAk/07fcyBECU6eaL9IkErAe2T5QF23Um1M6av/QN4hx
hR9sFVo3kuZ6ePmI5enrkQ+PL61v+Hvm+qgd9lesFOik7dZYjhFluSm59TBogi53
sl5mz6p0C/DQ9q8ow0/Ydo0IloNi270zVmHgLD+dRPYfyzEWRIgeNt3Udyl0OSjz
0IB5kt/YG8B6rJ0nSNYTY3uxSc4qIPSDjMi8oKcj6mnQLyyhKiHSRfFedMJE4tOc
l4SquBS/ChB4MCrH5fEzufL6APc1XoaG9Onqe3gw9aNVoDyznkebIoIFT/XRm2ZZ
Mcad/pk4SmTIMGEkt8WEr0ELSqMPzoL+WPMLZV9eCPXcbGe26ng8q0DtOhaPKyia
TxGwN/MjYs0JlTVqn+2GTKr9cZYP58VjCYjrYGm6tB30wNAmUnazP/ksRTWMm+6d
5EMYuIDGZ9+cAqs3fEhBSaCn4baCUW6Y5/Qll2Zkxb9w38qPdRg7DN5BEoAiG77w
ZVnNdgJfm2B97UfgXamKgt+ZBiy1HjtWlS7UdPCMDyFc1C6A18BuuiXyA0s8/JAj
fi48MC5Y23svAGnx3ud6RN+yKVQHT7m/0acjup8ARQIyl01Ro3AuP9+ioTpJHB2D
MQWtjifFwN3Xx9Tmalt7fyTrjCb+K+ZILt00VGBe/rqqpTdj/UBtxsTaBKaAxgnj
1efIgKL72qUVAxpZGkDjHOQ4iw0mER72NLVYEOHE53OP9919bCfyMj5WxoUyVG/h
X/5p8slioaeMw4MqR2nYk8cC4vPB25qHan8buZdu9cqR/oinbCH3OGnXJNng/9lZ
f8MV+tURG5Bk/zD2XRLOXWUPi0owKV+uxojjVZg9dmYY4ysiG8bj/74QF+/deaij
SUX//Yp+rf6x8ANW0ogxxlUaF9BuU14FZI93C8Zx4wiJkwZRaODkCY7CiyIKdvpg
vT1GNkYOIn8nvSt1VQXZ2bjBbLxUfYtbE0C7ov6HaKhETVuY9rRxc3HYnlVHulZv
+EWtDa/LmvzaFZ3+T3MZijsWKfZCe6DvbMBAogIAHk427lA1TQMHXastgh8qxUw1
TQn46PZXCc7Ik1T2J2zm5DVDzjDdlJEJgDVrjvU+kMDPqNJ37xGARUG0ftFFNThf
82msuaz8h/RSqQf75hE92E7ejzNf6IB66RN+BOPJt6+6qhvvep5i7Bmrcox2QpNb
3ulSj9G2hLBYeRg4iaBqABhd5mQf43XEcQ1AcKC09qlitbsE3rtQpVuphGxXN/0B
Sc6YW6lFbSBmqM2BsjSfWL5NvT1BVmVZ+RnYYMNo8w4c8hbFDYYlbMblfcNYl5WW
yCwenOj5K4GND7PVLeJmViH+Qk+kPsaR4Akhu3+SG9PeisrozMo9zqhhHUCpiZYZ
eqkM+fvF1VrN0EtCd/NrfQ470BDRT7YUvNGeEYiySXAvJyHddwbEiZ8RcTaD5dxL
6uRKOPs+xSTN4VILDpBhaxVCtyeE8CxSUh5db09oQ3FAlIYDTr63qU6OSPJTDs7x
2UnzyOSURo4mPPI2F2EZwYMCiP06aBzrpH6S2j/APNaA0UVv7Is/fNZEIEqhKQM6
W+t/d3yVok3r/h+FdEOfINBGBPuTK8fIoB/z9/bzBenjgvnD48jgfBx3A4bFHpLH
BNoe6HidF5rArQi+hasOeEse3wVvI24IbBVymIgIR8DQJcTQXHEIAJWWKyKY9vFF
HmLCww0wENK1wB+i/Tj28HwNg7/L36qNQZRjVPKLpH7qrFcwem3a9AehByuL1DBe
eYT173AmC5oi+t3+CfSeuip9ins0nAnkmSEen7q58Ded2rU2l+2MPbXltzVdUeCW
gL31iDuvW1WXvpNxS26CC1XcxEoFezzZHyFCjYuGHHLLVrSIR3qgsDAF7UQx0DJR
oUsE+maIwLJ6IdHX/1dT5HttuUEFDHQx8fZ3SMcZv1LEhsy+S3AAwGAK0Kvca39B
b/XQ4GAU/kj6sqUDveDWVkmPN0sFXEIKH1E9S+8twND4Zf27dktKmYO938iUGRth
Q3IOIvmuQZVWdq8h92i4cYPQ4iyaGWlq0xVuRl2x5vg9jELZPuhxvcYZ2LfWEhSf
RkWXT1A9sjil8z+I5LDmSpcZp948vEwwTxeDpEWLmqwt+Y5EiiFWT1M9PyejHeql
mVabj55Hm/Sr/6Ih/Uxt1QfMbyinNOxuFRb+ZclTawWvttBgTV8Zm+DNOjU7paG5
EHvQU5Ym4SxlavOfwoLa3hZzcwVVy6WE4jswMfsScJMqG0fzFnsVaxkvmoHcmmqp
cXup6z809mbSeZEeMPTMkmjotbjinuTuXxe9CpN5OyzJEef8FE8IywFmVYKerHOB
IPf8yUy3POxHaILox/7yjqx2QY/OcuCrK1JlXGz1niG82yi0k34kxxG6Ifjiu40+
bc3NHH8ndjFDqhewsGGxwQms7YHBReSsoD4XbcLKcratZgkWiri7AsqWvSFxBBBD
g+9tejTXZz5p3dMpJ44jAGf+ETFCpAIoD05o7Tiyy9V6j+hFv/D/j5L5TuWQPXjR
TnEunkaBoX/okC6HLdV98UHjowW2B34J31pWuvuNW7v5Web5zrb0sBc0twdwmbxw
30lkm0B0A7L0V82nH+VWUlWoatJE9yEUmLS6vmtYIczEeOQBsDTrlmR1jSIemNR/
VzlCTUsB2xvwPoXGZ/oD3KyDjIXLZeL2FihqQ7Zp9fBNkWl7wa2mPlZtc+eD2TPh
aQJf+pqudLCtJZ7mEwYepvFwIiPcvNC2uyNowkvW1hj8bdnk6PFe/YgAjmNopB19
nT8bVZ01+9SSk5dB4IjCxbfa8fF8SPBSd0UyOTlgw4jrURc6BycW3ZPvMxW9Mjly
GSHUkukn0zJiv8/m+wtwZDUdbm3xVC4Ba0aDOtYlJUzoPHsFjHtaJKRQESwanF4L
vB21NOtDiHgPxY0uhQoXIwAI/+yyr4FVSusnW4wncLRviffOM+Knsjui8gr5khNJ
cw3yJCVulLKQWuTe0DFqsUk7gclTyUbv3XL4dvIGcUr9hbt1jwXj/iPRTOgXXHav
aHQoiikUyLQOmtL1+30W644ceh0jPaB2GfJdFAYKkHDNpqwaDsdApiJZ64ZfDgeU
jUN+4Szj+tV6npQ5WFKWpAp09ZZNVGNXegcLe68/ESipJLKLDUEGjguwhx9WDJvM
mJEpGkqeC4uv4xqtJxzAkqBSSQo2ftJmWSfYXLsB+IjFAI73QptIUWWXI1kRmobU
FOhIMSNpIdmwUdS4raeZqEyOS1gtqajnHQxO/PH0+wtne//e98bKEYwWlafNkkVc
JEXtS+ceyWyCRBR4OuCUU4NbpmeuOQZEhb+wp7wnPnnq8v3t1La9qkWLP+Blnf4T
toJwiIsT/D1ZeD/GLEqzr7yYqE9lUnS/UXiGKgQ9pwP8SLCdIvbBubig9li2x/Gv
YC9RqP6Bq6UQrgA2nVil3QHasvVa6cwFFcm34n8drqhrxezTW4K+eQReFWFxMUcG
H84qVQGFcBcOHrFkJXUoKbqraxEDP7alTGPMJwh1UFrXJDI9gP6Glcf9YXGl6y/i
TW38vzlyYye1xI1ELkP0jR4fa1CU7GK/aWczPRkiRGQGjCE7/Z9c1gN2ZQaH0PEu
g4vK0F8X/pPc/9uiwGqxQMmMSmzzrT8cF1oSUImqY+CxJtycTiS7pDRmIOEyC2tC
A6OGfQj/gbH0yQOuTGwkZkwM40Ht+TEQUInMewiOFxd4hd+6DiM2Ifr9ZKIqdKqo
Tn6Y+u9faZKJ/KduF6/BFLUkH/OQdc8O/S/9FFJzApS5BEmlZH8ks8ukO8CQVkUB
BJC92ALC3I65sr9Tr0tfb5kSZicLcm4ldzAa+rcgsEGeepG793OEgpucrbhrWWxh
Fg4y6Vguemvrf9Hrk7WSm2qIBLOB45i+q6Ce4IwvCCx64C6zlCHRsRfzt2/zJ5Wd
WE07Ls6Oti0wCWYbP2FaJYED2f2+5XYs8YXtDg2xVe/5BX8Ka+bO82klCgBoGEba
I4+R3ybJnV/d0uuxeFboLdmoAj16W9InzBPlC6ESArzCfr7Yfwa7KCYaHq1j6LQt
aObmu2YTFkXaYRx9HTFII2G9SKe3fujZr5sQuxunP13+JhoCfa6Sq5Tx/89aMtZc
4sZGAb1ec3b5lMmSGGeX+e17eACRKHNSU9/X21OCZbLtA10ETmqjqnPGY3uQ8oN3
7Rc+D0A/tlrHuACwfeEPpHEiSwCf1OBfcl9O3lCfdRirPr9aX4Po2Am4i5yhI0o3
PhcyZ79+KdTBbxQQckQEuMLMO4NEdcjU5b23v55ZSwNE9W7sq7kHh7nlzrT9u3HZ
yE6dmMZJbr47IXSaNbae4BkFkYFNbdWcv1cGXj6/2PaOzI+PBzDr9zhl6cRAc+H6
3M0yLBF53bECM0wYG7LGyyGF+fk2YgG1lBWKLBOGYOZ9IWtMPj5sdvZQHfLgtpN5
MiR6KWxEiJ2Klk3sOAMXg5IiAaSXRevSR31XeHjkoD8jIW37pCbCFQyYXDXOqIQP
LiwmVVfcrB0et8Xe/wdgjoYY2qAlBwQ/s6JxQZabbQLlExokg9Ey4Hf0HOpKDjt2
YRbRCcRhJLgQ4NDD0LlvzdVsO6924krWa9NLjHtC4sI2v1ABI5t43inXeW+HmZJW
CnzLcnhc54B3IgtYgAhaBeyjAiIX8VU92iGQ4kcl8tF3zRUxq26Na3E6SmWDYfyG
tHYK7m3xTf7BNTkOwrUa2zRRg27ilj6u72QZIFjuYXZpGIDj+Og1PRFaRnf4MDGT
QitzzN0TCnaMV/0/ijQrSAZqZIKtbwNIABnJem2G6VbjiNZ+EPPcqWOn7/CMd2yw
hpoV4yg4hbk3U08hC7+eibmOeAfEVlBQ99N41NBdm9F3r3gUZeYV5HvEzxZhsHn/
g053fXWf14++TrWevQUqrJ0rNTwK/rmKYWcksOpfb53/61Q9Pmkcw3ktHeKPVDQY
HUdqRwcoE0ag2/w7gGeNIdjRxRTAt6X9+NHmPK0uVrVWEXIYE5rKKbB/AipMzAkp
lqpWwaj1YLNzaHzzP6DnYHs1x3m6LZGsYj23p4Mb5BS6zxQg7ztwQEj+jnydK9IC
UOErlIz6UY0vG5aErQpaZHKkx9xLp9h9Q/KSqOY65KmKGyZ70qHmnbkHP9gQ5I1u
9RQo97HubvCK6uk2eJsDv0ZZDC8SvHj3v7l4jhYr0i1nehInTf/9FesLLleS09U4
CybMmrLiwOPE79wfr3EiCGutb8m/m773d5wEHRdvv4Z8UtUUfsIGeHd5MUDUkVeG
pA260gmmGX2nz9dykl89JmLnors3JgN2+XeBdxl24G7+GWk2I2j5F29z1lzQcUV8
eiKj9njGw6fK6jiGXNz85VkVwk6xwuEjrtB2baymkVvp043JPpRazRlt4g/uZmAB
IR+hT3EnjUkjSt4dQHKrY/3qOtL8fjui2K3Qp9IclAoANW0oN+VM2oyzKb9plYkM
MClOHL4zQcHvUwPA2xnXavudoj/GuafMtonystWgEcgghljs+q3f1CsoBNUw3rfH
9FuWzPbuu0cNSkRju122vC5FYLG2JR0MVCOJF5dsoU8oU5GU7O0s5WKZioFQJoU0
Dg/aeynDooKGrXS2hu1Pwy2fgvHw6HiHC9fhbxqtOTdRlJ54ajW1IILeQ2yxfilr
NtX6/hqsxy0VN9f9RrXUvLyIZTMiqeaFkQuoP5qLUG7EyxP6VlkIwP9TMhwImge1
W1SCLOJsWTn9TlkSuq0G+iGYCTvb9aaFTk5AwP8+uE0rpcI32+/X5aUUYTiCqhWJ
bEJmZ7gbJVysHzFZismvsoe1Jd/4s0cFNm0hn+JSBsKZXUGgd+4EqR0zCDXPan83
M84Joo1cOZr2FLOLgwLVGo+PZU1dBV2BrkztWZUlR+ZRLSEVYEnyVsAUDU1XKaEN
F0RrMK1dApE+qV9WyfVjviJZnandNW1nWnccbSFxbob6ByyiJVtvHIsD5ZfeFSwU
fwjzAYpUzOAg+N4hfaM5esX5QmMR7WBBiaplRcqnfXs5Fkk5HIoXeR4k6QOeQ8ab
otQE+5UJkKxJYsQLvOd9UdDaUF58QOPAvYREmMT8jNoRXuY+za/tR16KSz38YApi
ij5ezudizfKc05YwDNPTMWp9VjSGiecT5S6VabS6jyI03HHFBhXNxdQfQIq0X+ou
qclAJEVXJujXDBUwa6m5heUkRnzXBgNcPZFyrINW+/b2ENk0jsI0imuT3aOyu4cv
/ZbRAKfRWUBNK6dOJE6t2oO8b8cyz5huaycItUpGSGNtMWBWbMuTThZvxgXf/Oba
1zXXXAVkxrGoe4IPkGtyRZlhzwt6mWDfzF/gMmtcnLSFav9RTWDwTzCY1tPMd19L
vAY/aQwOrKXm+wL1nCkjMJrVml1YvfIHNtQ1cdXgjv9FwxLv97U+Z8bEocVc7gVn
42iXlOY3rdmDGkykwuZRwz8sduo7Y2H4xqvNYiXFrmERsL9Vr4wBAOSS/RvB9KMX
PEyC5KdeifrAI0Ebz+GrosGSnqQ/NhsnZq4wFyOcpWopgP1rKK/pOVUurzqCbNg9
IddavYNMdf1kGE4kdFMCTxRgwljdxyBcNudKYTMV2yvz4S9S9dWC+RkIfNoo+NTG
l6WEvQfdffL5IxLvcNZW/UBPRFcdJsgSALOjJPNS8NxTR+fGkgcDSqpfu3jlZdcF
uhfHn2plaXDIsTAZdKLrh4SI2NwblAWCo335Niliu7UheYtBrlf87pg2y/2ryWYL
8h2O23VgR2K8dHAP7XtBmvH1Al8G8WqfkYawLfEfByNSmY7E3zdKvHAOj601UiRK
2juy5Wy/tLS+ysZNl2aMbo/na/KcNTy5QkkhPk/kQiXho1o6Yv7qMIzujCDuzqwb
e9U7nIdBaPpDw9woj8HGVgDi33rIDodXp+plhHxEtxL1Qp1n3kZx5urtirgkzcX1
ot9r1b9dXyffmRLqUc9GD5GNEUYC3NEz3RVAtr1KCc+OH418P+UesguSkVAvDG7r
TGBO+nRavBwy+2AdfF67Qo0RoIRiqoRYgko0PfO3vgPf5TYps5gLgCJlRD0B5pIk
Rv4gpWIEbLTRvjICXKlkHR2ynMyZcz1ij+Un8kM/9TdBrNf2LkZWn9pK2ndWU3kD
lm/QCu+P9OiHe9wa5stsF9JDsuNBkRnRc2gNQrWg18Zcmx++847MwnjW2x5FeHZm
Xrs2jxAMdYSMvWYtYIiKon6irZ+ZYPx7rrdp86ToK6uQkFpUqkkMqzNt7EaITOyh
TjF419A3RJsnuG4OHtADTzWemzX2aBvEKpgZslLhLZ1fq2y0NSvMjMMQkzjeSrO+
peppgqNJU60f8o9+UgB687bc/ooyKZwnmx9n1sx7iU5xT5jwC3mNAUMECI4StBnM
E0WUbgDvXmkIXTh/DJ+NwkmE3awJXBCS4E1/8YcZPVS62zKImvtIR8ttJDDb+tVL
DLgymuYyRRiOo6bMnf+Q9g2z/p6sqqFU0hoGjALzY1Tm6Rukjni9eYAcch779rR7
LvxbQaWRw+TqYaSwHOU1CMAhPtf6k6fCIwfypXjkGidOLT2Qxmjdp+RiDCE+Cgm5
4E1Kly5stUIXSckyX/200Hdh3UQl7Rbz42n2kWkAtTSOPILA7FiXRKN01V2zbaWu
rzMjqBaGn8OG/WAGJsCjmxNI+1mZysyBFWya+A+nKY84UtqWVLNynma4kKi8xJif
nPn8FsNA3h5TZeb5wS9id6wCSadx2cFFaWUfgn8jfXHF2pHqKbbzryc0v0HMZYlr
i9gcKuoXLUmCP1GR2VYM+6qHsNHvsPJIHyqJJrAAgrkyOfP6CayYvu+xcRxI5rs0
2CCTgUKXU5GJRyUqODnqLysiiJzcrUCKvB2bxQ/7faGd71mT/PG95/1ll6YKNEjD
42GX5kn+TR0cDQgGubDvvEeBevwlkecOErkBCTdosrPP/noel7gEw45bl4dwD7TW
2pSmJq2+bGKLa9JZGvAl1nxk5QE0d3tqRNsZ0jwCVdgwF1Gu3G/8kK6ID53lrOii
ZQSMqCOURHo34cWWKrcheD6ei21zae3ihfXeIi/fYS9OSngL8M/aGNGebMUr19Lf
7HrK6QzWh74I3RMQkSlzfXYx+SExqLI1p1yJKqngod55lF22kpBCigrhQTgRElyP
fr3IJUrdBUmP5VOR/w6erIE/5Z1b2/N8Ec2+SXVGHTJ95vBev2H6VLB01bpC0Esw
P/BWzHRGwWN72jaBmSbte+R6Y6gQEBUusHvDWb9qYpCfY4CYCk8TDQSHi8dU3mUr
nz173094LPdQpKVS6y/rHEgm0s2MG8GBuTsGOyZElzYBRMFcUMtqXGLGoquLrBsR
44KTb6mZbMII2LRt0sE4ZihNFO7tmdfs7nQTGlEV5bvfgnkALXkhrtwFXJvbAIrD
Y5ahSr/RNmRgvfoBWaOyx61f/g+PN9HnAAabFEbuu3hi9vexdoPEPvbAYgrVr8Hb
UIAne73impAn1gGHMYOgmq8rLC3yZKzZExqg7to8jzBWKqSe2ptk9b4e9ht+e/2n
WkhjuGmZiexYOU7sWEu0AXhNniwVlzEG1Y/+TH7mtZq3TGMbTH6CFdcVY4602hkY
0bsNxpTClR0PyQUPmVRrzr7t4goQ+O/ln2aKvBRB+Edw9VkI18XBdxn12Da/T6na
DU2ApobXuJy6nemMuESckEP+KAqTG3/kg6Adxz8CnSd3zv8XA5Xtn/bG7vI6vXR7
W8o896nkvL7dS2uHBpejv4RE2EdSHWi/jH1lfp/Oneijnt0G4H1DQHAjwqHHalUu
KRzmQQrbuJXPPrBR9dmi3dCC8jbUaG5u4M+dQEbaTeSIA8s6aEDdMdERWRoJyVvS
HFwsU37efSBKjeCMV+Et4Mp43sqvHVuB9N1Z+9D8zMxh9Ip0JYWRdTh7G/qkObY5
O5CWNn0g2Aml622tcvajKAFAq5/9RV8c8+rAwvSR2UzXkqEjIO1CvAX5hbncAaW2
8wf4yivGR61ljIOZaY38WnrtDuWAmDFjVWTT+G9GeL2viXanb5Ei/B9P5yYH3YFQ
naXylf1GlKMsvPy0jiGWyIU8QBFz7e2kfdcJORWBe6Xa5s7wiCVjDairRwAk5Sdc
cCJv0HYQQb3RIYDX2tmzjkTkB7GU/fk8+quZrrsysAkcMIpM/DJb/EKpWTN/AvoD
gDpEf1gRcfTmYcURb5LTzefL5D8jk4t6dCam5E1zx/JLy/dGf0DWviZfvxyFCWVc
gz0HHF3Uf4UIjhALKu3jJazjqKsmcai67h3kHTaDpNdxYbUpPEfyQpOdSxmebeKU
3Tkt5Ge/6Y+TEl4xjSjUFZrmmATzH1wFdVX7zItKly2o1VWCd6HJdIusLskaS5V5
llAtu0WHc2ZjM4o6Vh3olO2D3zdcQXLerFeiXn/XvavPc3wkoq5mS34ukz+EZpwq
/MlcWNvZlT+U/NV+8TQgpxMlxYu8C5wPs2EKP7gB9pxb3QN3KAhoyiHSZ4sFCxKT
FHPsShH0cJQKFgIWx7UpJUrdQEgQC60OVgGDke3Zlmw/Yzg04aX5bu6Ks9lpKfP/
1W2kWW1c62sPzqK+KMK9a9ssPPdA8+D+Q5e9wOwO1nmVJRTme6+zgSVdbQ8ou48z
I70T4ZmZyCHfo8JbnCUni9ZXkNqJrvYRK5/XbRi5/UynWZc10XHEKElwaWpgVfqv
ZaS7DD3Rj52k1l5d7l/HGkeZfhkXFK90hmKQx9nzxj9gPnFi8n0Y7+2wSCW96ehv
GNdwqEp7QqKePCGjJkgQ3xbVujWNgMb39eh9YgQUzYnfvU3Cd0jyW5SvYJcYBeYA
GfXkRdnDFdSQiuR4NKNjYVUodvAg05eYwuXhK0vKQfXlmgVMWth3hWFCZY2ohTLs
4eHNmb2MtEUIv5n/akgI8LeoibgHB6+GnSQLjvU13OdWHgalrfycz2pCyGKTS4TA
uSNHZ0c8ugU09vOlgYFYisTgaqYSSVz+E7Q9VPinq+1yHObChCh0i/t8ZXAAHLAz
rN8VX0Aqjz8ENOCdZQIQ/cJrde4270kV+exnXAdLo43Azcbh1oJYeEyeJG9Ch2O8
7EYWVYsrlZKG63+n6h+f45qJiAIdobbDtHsHxF6iAx6biT91OybSttj7QK12Dlg/
kHlmLmX5H3j6hlA7EJmTpKGgklZ9auUuqciDZIdqaiDeLNMFpJH29K+cJuadkl5o
YgorAovipyZ1mkNUzmPEmh/ghQvXYg63Uzq7kxjo4k0LFCmQCHIVjxsk75VBty3a
cIq3BRu9UxVmjXkamI/HxFaHS35aEAPIEkIYP8YJWrqcTE22WD7akhAz184qh/6O
e/3kNC+//nrSrAoc+iWXFGE5kcEYb5ZvJgPfUxUYclXHBr1vmDbNQa+usuEr3q7H
BTT7hE4/nkps30UvPbubSi0qCnGcLljecd3XWZ6aH3VAUz8QH5p9G4TZ0H/PGehv
XXCEhbBNBzeslJjxbJLh0024Ys5FPuPTOjbAC6EMHCeSSIMUFA3nC+/rdNPEA5b4
SgSvGnQldmjI+khPxLfJzm5c1N0c35uJN/l2EA6Z9qwB3M/KCN31CBVHM0TVMtnr
Mp914DVAmWPxOYKT8UrZr2pt+XAPBjyfWDxkuvJMZYPMIOdMQEJDUZCFr1a2Df+m
4EHa2PeWNFBx13VtcBELSPateuxxMlPUHkEdLqGzqcJHoM+XBmiOENlYAcZTIEVA
vA8JpoOIHHxsM6rNqK8Dlf4YDNiUZIxV9dc5jsVgn73G/E6D4AoIsJWn9nsbS3/C
qc24z6G7vFJlmn/LtxUQ6E2FkW7QXjMVVsXFCoGPUznkk0eXL8HYjJ7y7gj++J6Q
QTRDQz9YbHzGlhjTYd8mHM0AHNkhb4tEyplFFK66poE7gMiAf+VnDIkVaCRW5EhS
AaI7pKisant4xpI/gqffTIv//VgxL33kcjzIZhz+A8KEKhwrplESRZbpRW16UX8N
h9bcu2zJP07NsvpD6g93B0NsuaodqR+vxtQm1APylxo6I6kMouDY8YqHVAFMoqWe
1M2gt1kDehN6G0nUgQwH5Jc8BwCnNGIR0nE0snytx7N068ItkyQtVvf7QMg5lLAS
3iRvAsyuVg4obfDP16egB9PYgf4EKIhzXH4SQ9MmpEn28+GCqe2FOf4uGlSPyOHm
dIXKj6ysIoEQbbuO+99Wks9nlPm0PpO0MLHYTpO4FRO4tCcAo08ggxSrm2kDXWx3
OpNmbT0OV1xSmgcOzZ900vhKA4mXXxJYAzTlNfWHw8HPnRXPPw/5CA6sXVPTGd1L
D4s3VXYoNZYlwBXz4LmwqYNnohC9vN3la1vIbqzYaXXYMCBzQe0NOsjo0eW3RP/A
umEXJzWt3eAhOy9DbynRWQ4eKBUDmL90htKQvk9tyaKBv/lUa3SzOMC7UZjfdI4M
hQwSMvM3p6k/ltaJQjHM3GkfYhba3+MUhpP+BTnk1n1i8ACnaFVm95HtJNJGLtcY
rNvU5ncmT3Vviqky/jlEFsWvrU9IV1i4Mq/OLDM7VlJE1rJ/XFa+suOIrGhjhj+v
SV+I5ErsjUHtHCiyW7vq8N8kdVZwKHSD3UuJUH20JnaVNjVsbWI6Sr9JiIONzm+7
SglM9Now1BAFJ+u3gvF53/n9DFIDEGD6SVY0oH3DSvP8mFdnXgR3g4NZzkqvLDA1
7dKUOP5xK+mqoxFrgt6/F+LJz1gD2n9Vgj9xNT98tkIMrOxzLf1cl0gp3oSGFGuJ
GoPLU+EN94NXJS60VZjSS7pwdmzAos2eN9p5TWpgCju/pDLpbJY61d5USabYAQT2
AlUUEEE3TvnhyLCdpGtPWcJLkqyc+tE1qrdDVoo5ETlDKeVPdbseZm68PpzKoXAJ
xA9e+QQZgw2bjMjVHmBdih1Duh7EmoOZ514FJlbxD4ARU1KNyZEzCybzsdtNZ0oX
gambrgArFlkzNZvtwQJfzP9A4iSGlzUbCWv0hqyYxY4m1VWi4VQvqSSvg+9R/6fD
/XwfkQ/p2rUmHkiLLRGy8cl8pKEMMS/0weNpsDP8x6I71rdvi04MksVRB0Dvuafz
7LhDg7MkMR/bYGn4gXEs0u21Lx+H2fceaJTo3QxJGu60Qz5CqzK0hQGCal7ShMZm
qt0e0yM4cQaqAIikdI8sCHWiN4DImFWmEesMHkav6OhpUer8+A/QAiZc4sQqL4Jx
kLKnalS06OqgiBu9aiZHiLuVvW4/Dmr36Rgk9MId5CpqC2ctAmitKvEqEvFSwN1x
oaC7BBR+1YGIQCNsnQd5EQU/3IyvPONQ8E4QTH+PhACp4qL4lbsPJ9qZ34yFleY1
UH2VDORttRHOhHppFqFN4htzn+Q5huk0UB+X95/DilywWeVzPEWZisS+VbP8Xm1n
44Eo0u94nILb6RN6AeCKQc3v+cEDaSYUw6/exjNJIDFpTez4iTUemJb+rcK/C0b0
PM6jPZKpjAK+EfCL4JytCY5troQi+iwL7N1TCQbjFg7bNLMgEvfp/PMyaJHJZbT3
MdjM4hAsz/5l5rvqYeVvap+MA0E6L/t/30hZgy77tZrt32gVDvE2s6hqyxzAGs7c
fdyUxAQ57y8n/ylmxWQScGJofxhiuDEk9A67QdsY13UXtWrRcL4KfkXOMFDQKy2O
q3lGWv7tCpgbgLL5E2jFZ68aTeW2gVTkQ2XyjablIlkar//HYZGKL9FUcH/ThU/V
KWJ0/iD8n37iU9UDmTB+qOXK+kt9defCc+sXkVXnMibfO6ZOYJnc5HFO/FU33Vzv
IrM1ojtAHIdx5GEYH4JtARVf1TQdsYAyuKQzdeObA1l9olX5V4PZJ4quaWiYPIhD
pEZGQSst0nZ1L7d0n5IOwYAfmhxddJ/TRyTzj6NYLWIJtBIIhMOzYiGJEouD5YqS
vbYrd7ZhsYi33K1avrsexBqTqCowL1rsgKGE3ayXSdI5Vaf0bB9P3+gtq41i6Q//
o9+SXByTAHeIlrnm0idFKfE+y7AxZslKajGenmiJC04zjX6Tk4O6HcPMQvF5I1Vf
YYASkrwRTl0ex5InKlZMGMRrwKpWpVECuCStTO+VugOm5a0gV5JGMBy90UEiC3G9
y4Jqgzx5b4/mvjnssrUvVsKBPG7DVP9842mYfnx1aktHvVAGQEhEx7I9wWENF8v5
N6kPocuFz/GjRQ0Zq0D0o0t0zLA6viAR94q3rRkEcwUA4Pes1ZziVy4o+IEY+Eph
fkoDXlKzd+bm58yx2Iyr4iUO1H/maN2xv8ZRLPry24x6xQUvORtZHVRIpnZnkGTC
VGTIF1GyGL3tP6mG3cWdC+F1fSU1KXuqu96OyXDvIuj+X05FtA10UW0InnuDwRu+
HXEpWMKJArFysSFx0oUeE9eL4aYIw7xEszJIsEe+kT5RftIwRosQ2WvoOSRAWLsj
SO1Q1Kmg90TvbcMjOAzTC5NYXgFEYy5l7CTn2QCAfKon2CWS7qFn2Iy04ksAYIBe
a32djQgwud0BZKRbeZulnVSkF/itqqrNJqbmpGKKqJE3Bxh4a0Q81t3FViv81m8T
wP7WB02EepEJHi7vXd32afVUkwyiqU95Jr0n9wxrMfrPKl7dJcoKTpFbFlBFSyLU
a5u0w62/r1ozINIqoGJMYQEE9KTUjRM94Hpumg8dHzKwvuGXhvLoHcdwF7tn8W7d
wBH5JWS/0PYMmLjYSIQqKculKxUZBam6zeGOXTzmVTi0/UdJiQrLG+2nQRLoGpOU
91cxGPFbn3vRf4ywyhxz+Q2/Pu1Dgox/aglqT8kJTdVrdLWurgSlsmYx06FYh//v
nXAdhZ/wudQsHU/abQZdTGGDMDdHBs6p6lU17rhBI+VNyIdblF897YU26Ivm7Mz5
aferGUbLvGGTsnlM7oA42QpisIDF0RX3+eFEQBq5xzMg9lhpz3bqNAgSYkNACOpJ
fwwtYEyonylLwsJ04K8G9OCXl+kwzLmomypsw+NLUD9hV++BIOkOIW8yKFNkfn9S
BxkisQ7aSzzo/LoMaWAuMBl/KQLiWK5K8GRu//Yd3E8fIUxIA2FWaaoqnwpTlmFB
Q0b8yc6gHpS2+7ZpEDaBOwelt/ByhNz5UXeez81W6EPiu3xDbo+fJVqBZ9lOfbj6
F5icOMwW+oqqtWTply3UXQtnEHYJnWpJxSc7IyH6WUa+XyFtNpVNcMWvEefWPrGh
OBv+NUgGEVflcqrRwhhRmDBFhfPXTToXv1N08fpTRePe4Q3K0Efy0dt1c0V+tbdd
SebPdtDxrbsJcp49fsK0podiwUtKI+HWbVfECs8GZBq0B1tUgz4m0dSv5bmAJ4cv
8ShaEJReoGb7S7j9ZdYxciicjQy+UCKJRlg4u+HrEtM7TlCMpuH2gapFAT9X9Bdt
6rOACP6XqCn7UDbfBn5jKWbtLerkGc86EI3ln79yAeyAt1WYNgLXdOdeKr9lIwkq
gMhkeA0h1hkOjVASn5ZHflC1cyhl+cBr7a4JjKEbWAxVClnCU9uLyZnoY170ySw7
N+f4Avbd0bxCIcwla13imSSRTzuG7L3iP76FbpWOzBBpWzjFne0JYCeFVnxpTUu6
fW5bS/0ebfrLIGYJ/EWYaI9ZQ8LktfajMs4Q8dsPgdDoYZZDR0SMd0A0ANdaqxFq
fdhp6w7/u4Y1Q+wYoz1mVofHQp6Ugq9xvGuiGWSfvq3BXjwVdm1eCABDMsaR+BFH
JkHS0rZXA+T+LlS3mLJjrd9+0LHOVUmBrH+UGSrkESNfRTwPGZaLgXlSQx2W5qZg
ABxQpf4SkojNe/U9KL+YbgkNIa/vl551gByJHuchia99VaJVYeVhNI4nyAc88zc3
P2+ym2C8zYuFbLa13PDF3fc0ZORlvHlQQ33crQDTF88DqJcjxfgovCBqy/8+4BsC
1gP21te9DJhpS17Vq5GbPasmjSfrJcd+O+k781oHfVLm+TUu+aI5/YBfoLwagNve
XUzL8huTKI0wUAQBvv+32dmirTboCtXy7/MFJklebtXscSSdAkK4MrjzDtsUf9X2
sQIenKq25aFXgMHXKv/278I180TBcJsBDHsuj7dRWDQfG95wEQzx/lOIBR5bshSn
LuAcMtG/oEFLGBczdr9xAgtJ330KDcV3s1zAYtwEiA1pEZEv5w82sGo5U4GnA62F
d5Ugy0Y5iunIoVnJiz8vjI3589esNHZ8N2Pd4g97FciBYBU1CkUwd4aKy2K069+e
F1BNfqL0hP4mP2LGu0pplf0xc9o9Mc+DnOaXF3CWI36QGkB+eWGMjMJi6Ibzg71q
JAUW0hNqA8IJtjXQ/1PVYc2CX3gcskqITHzRDHHqNzL/I9Zp3/+9jmIFHxWl3vv+
PiFcdF/jUK6unGb+a0IsGjI4ds3UHUVQJXFV9IKIMGiWXzuvQVeOrq/jrbTyEanH
QqTTUiz02+1zGrq+g/6kog8asLxBvvmEVwFqV4khGF9/rkSJJFbINGEPCKF2TsFM
N9BPwZ12cwJ7tLZKwmxK7cKPMfPhtU+vTa5VABblR1DW87pF9RZy5zGnnhGD83go
LFZoex3oS+2UVQXTXVQrkrtzHPbSI7T35siC14umwFStFWuWinLBVJ0Hgw4wFEvK
D6B/fyVU5d0Q0qZU4bbT0zXUBJnvUG3dddJ1sRiTvP2sk0n+nohcSJIto3Tm8YCv
1zrHxd1yESNCptKIaul6x59XSPRypXyzRWkvnzO3X84CABOe66FUgpUrQLMqUyfD
TmRt6NnejQMcnry0BsciZNK9ZIk3HhifNxNaH6vi0XBejl3s1lai7ZJ3VDzz+CNW
56GWIlDAz+4Ab59GTaOF8FXGGGYhF08Tw35o5jVM4l1dg/EAFGAH1TG2GPxSzjbl
SzU/f6knA+hJWvQRopMh3QY54y1mkV6I2d5dNGBYFReIeeKF47jQVlcsC2eFlQND
/1tddtCjJ1ObI2ylHZcRfhXKuzgexkee1G8IO4nETl9ZY8/AkrRN6Lc1TgIbOnJu
hnMKI+lOMsLL23MdSunJ7RBSkt2AhtoX0099vN/aKkrE4j08OyU7JGWwTwNu2MtC
HyAdy2/U0STrzSx2M0y3dGjPMk+JJ+lgSRaXTeAcJK0jvexLeQgqYbMQt+teTFld
r+qCpBHA5uRVeYFMl0MJZpbLtMTc2QxoQbAPkuox1y3Hm0ax21SnX1R6KsqE4NO3
edb3t2OxGpfr5emawBheTrVT5QOixl7Pk+RXQHaUjWcqD/YvgdGdvm2SFgQ7U82L
F5w6a2Whjce9H3OLZ8+up6kbJMYzFDNB4nkuTfTWml7sdeEeIPfwDhsZjx1i0Z0n
JsIJCm690hFnvI36342kQsuq+kd0IEcWwP3HJxRQEWLs0Dh3dqBBGZo7RP59D5Pt
898ccfOldwOJYKvztn/nIHAZY0jPPdEFKhSeSDzXN75yr/54KUrtVzE3II/kctu9
BUIyywa8XXF6OCjGx2N3mV5yFbOHDdDn0KB7St72dqUzDLj2qfMqvfJuXOocs/Nq
CNwlA9uKwPGhOQ1robPsu3tjvJjZFHwkegi+O/Wp8bmQzmkNX4uQzDFtM6B8xHlU
LE+CqSrKCN7HZaMIcADbFaQpsgIssPe4yNyDbdEU/Vag+0C8hQJG4q1JGbE4Om8D
KkOcp28S37k/eDpDQ31lwyB2QEBaaeGmiXOQ51hEn4kD4JRUwsY2LCOypRaRuGf3
bVrS1Sre0UdPxEZE722/6b8hlkGf1dmKldJyp2xXcGIq+qMuirSOxfAqaj9uhLoY
WVD//rUZL0wk6NNR445pyUw28IDSbOyQN0neX/pgaibeKUXDM3lnqMWoCmHTAlrB
tuuekAeIqLeEep0G94WYPURBZSiawdd30N4N4QNl2pVdpDjSR3C+T39U3LJjFmLW
1shxT52lS6X7pQ5LUsi+LplZzrA0A6tRLwS1Czts1FNvFS0QHyAqbitvwkGNPpjZ
4fuPAGkGej031I0o6MLMZudhBVaEOgBdlTQutRATl45+Hi+i7iO0TwPzlcvUacMa
SoxFacC+Q0L7ShyBNd3GxsvrydwRbQfZ1FR9wTMLvu0GxU5UbqbGSlWGvX35ctST
qFmkICouLMQLsIpwCDOJA/pXIfj73C7+h6rkRSJI1adn/1xF377V8tMWzD5daV/i
bveqxXwKIVodMn3SIOLUvpeYLBBvSpJx+rO61t1o7/KUwP5sy1bPIo1olgnX22qq
o0Q2xPiUYmSe7cvvuVJQZcKosf0vw/6t6G3XBnzrpvOcN7yopx26mw4Xkhnr4Ylb
MEg1bmKW/HKIx5azB04dQCEmlbU/qCR+btINmzeBtzH0AsCg53Q+neOjCuCM/6Nw
X1DpljQ/aEaBDTgPAAahD64wKu+oxy/jCQb9kzwukBx58+XmO1puG7wb54WDNanc
lclxATOQ5gtvewVkr2GaguwnPSg7l1c7b+IJkn2i6DjfWAC5si/th+J2WxB9YvJW
PHk0RtphP/1E1Ej+rOX7/AMtECHzfvsc4q9T1z3nuOBrD2Nmdvty38O+9KSW/VeG
ibD7NpBS9pIuXcJiCR0wCm22qpjjFqjnT3x79UP62q/rEjTm/AmQRYno6ScOttWQ
Bd8l6NDdNUAulC4pnSU26hiVyRKHH67uO5QtW1GEdDq3/gaDBLLBLX8PANE8vWFY
++qIsH9BZi78vdg57/uypLAaAgDPmHNQry6WboAVbEp+NSgZ4OXuePFxEXP9/iN+
yEkAPYU1VBrEp5R55LIGjmwP3ptvCZz0DGy+15o+RYzau3UpiKHq1aebADP2FvkJ
ziELonaSmo1YKv4YPhVf0EjAfUZ07XC7Ng+14okhx10QCItp/pXPr7uau+oxKVps
qVyAYQMyuVv8ZuLGHo3cKLr1J1/tCmEgWzLAjCKBmJzua7x7Cztn+SwEaNpKQiSt
LRnx8vj8UV8yOBzmxJrh7ML6kNXUCd6zEMiljN+N6/MNL76v1u+wMkpb5xec0vxM
H9xb2Cjvs/dJrYPOWt3dml4nRRmIcply2fxdCw1uPWqoiiNDRYZgZDeAmgb9OM2w
wk5JmJMCYwGpDH/V99XDU0aR74/A4r4ZLRKX3Rykq142qQraCysqq9dmaFD9ykTs
7DOO5oL1aSBjGZqqcpTMDel2zWVpdWoFVo/snbt9wuNWW5plbV0lVCyOKGcAVfzq
FkwhldlGp7twyU46i0KGEIh5anvaVJ2mNG13cezHlUEt5DReoAuXqh6Gn4InFfpv
59byR7/2cCL0R6MV7R3+kRZmFmyOGw6WFEo++XnlOEvxQlYF9qo47a+xwdmIy7AK
lpCM7kH/V/yrjEAomhur7EeUzG3cmWCSsQdMcqPUA9dkr2yPOJm0MtPOyl0Lbb9J
uN3h/lnHKsJt29d4+c3cOSw5YNmgc0U1AAmCkiTl/73vzIMx/02kZz7iZXDE1fxe
EeGEG5StwOG9AKvvaUlSWwl4ifBRUcZI3FmZ5v5cX53ORbOeauxisljEuwnZuV1M
MjiaU3clFxsJaXuZVOfbTKQYi2A0tWmDPYcwotU6ghrzVe0bNPFmbsfXQ4o2HDW5
Rgwb25ordPZ4Qc3R1Xhdk/1cxN/5CED0kjdeDPMyvDEI+l5amo5sKVevYYDxvn+q
aLi7uYkI9eLc+PEWgjfoANYO0RiiZLEVUKBEbWZGNsbhD6mGJHHfji4zlvCXZJAz
ZRtYLu3si/M1h+MesfdDUyvwtW3X3NXtXsMtCcprZx3zJi/wvT8F2CAnmPXRfHT6
swtSFHJmJb2XNxDlIR8TtCAlUkfd48J6XtHfaQ3Fl6pkwIHkqKPQNtWo2T/jwlFg
QcZgjV8Y+Pgq6g2u373b80emJVG+HQYiZcC0NsfcsHk6EHJn3LnYppcldFeK8X9x
uF3SjNTBfDZX6fZD7O3l/yDmiCB0jht6RpuCAzifE2sccjb0XbN4HtEdny7B8wHB
VFwA/XzBPWutDKUDRx6+q0sHOCotmrVQkJKDFnz4XohQe5zHIcW28zOrWpeJexoY
cUsYcffcCJC02eatfMyUCuinhk7KxqM3kmrlrAdx+bZIK4zw2GrSvn5yKqPpSzO+
AzJkK9/ACPcAqwahodWUVXr2tv4d9qzGEvLgteus7lpe7Jd0oC5EsCjqnqnHlKxh
nUkuRuyC1gU0NLxmkDsRnN62FTOgz1WggqvGgG7bTk7kU92x4dMJaYgVIGxI4xj9
4ojH2VfEi0QnHcLx3uoArMXmhYZCeIw0LTJPWARhWxdymT6sguL1oIr1DK1jzZ0W
k3ne5L+05GeQdKQESDyfYmeEpj+aYtregKO/3zFD/JskMoaS1Ilt7FEbOPbNqOyy
O2h72ualaugp8t+rx2dY8AZbJ/iJNPL9cClVg2ZEpKo0ONovTOudX8yytkAfP+wP
GuTTHBauwyTOZbMt6ooR4OVKONtgOd5QxdWxJk/V62a857EvU8ifb4IsTsy6TPhG
6z7RXp3uSZJWZuZVdu7V2dvvj9yDxZdm6btkXPeQnA3klAjXjMrfJ2BwYSBeHpGQ
7EjbmSqio2PzPqc0WyL1waMRb4G5m0WdKuvy8n3N7G72wB6p8lUCs2mDwgmMTeJo
gvVPHQ2H6lKDP4ll3IjlLeLnHOycwhhT2Yc5aWWSteizN5NHYpBxudIOmwrFC/bP
IOObEPCyflzivao/uysiBQIwY5MnAvKH377y/mj1X/cn7jsAvfk8WPJJlmTa4W98
i0ObaNM0NdkBaP0ptXn/UDvKf8uY+wq6sB73BS6Z2sZFIASd1n45vHCXScRwYUv9
xsjcvlP3eg21kUlEC9VIQjrq2KhqnueR8I5r10RFSltXkDUKELcTrkctw5uZXM/u
Lv1+0WC4jpjQl4GO4gXOHtTovWRoDDqHxYzSyopPooiHpctAaoAcf4IyEingX7TE
mF0zfIjoGHeDDd4ablgrhl8ZpRj7FIkF6h2ExvTME2kfIMQmSd0YLcq35Km2GysE
f7dxnGBYqvofazD9A4WQ9fLKt6ASvESLMhCTWoJ/FSmnGZ41k0T7wi6Yok8Np5rL
q47FmB6aXsQQkkXU7F1aHPusSv8ad2GDTOhtwlKvpah43MoXHO4yIrUYl6lO7j6X
c5XR302GLi3Ex/KqG2P5Ut1gEUc4cc+MOaTwveVbaVkDW19YZvoM2kpHEADrItiT
AdC5TZZfkFKnCQ+z4r+5q9KtAyiw4K4LJ9cR7KgpXeOvnwiXdRXsHXQnHXgBoMC3
e72adoU2pjvLY5DCpZqwd5E/my6sfX+TaswMeN7Brza2DhjY0EmovdmQ0NZg1EFH
gudoDREffOHclJ59vhEerS9OwcltgalyafJQQdh2qEXRFPytoQoFu6fNVQl+VCkj
XmKyt2fihGZRu7vLRJ4zs/Lz2A0ZwYpfhhDCmT32G1OwjDULAKRvfbgGbLkwz55x
ck5UNVWTIL7ippS7PFpM7Dv2Vp+GCdaFdLny6FQ3vZuMX/1XCCyRho/crpaDNDhk
DFnxksGkqtqRnGSOwbQwgIwGDSXi1CSyKQFkwSM+RNr1iSgW7s9MxXyJsL/o/Ua/
VoOeJHND5Y6Qcf9Atlu2h6Bsh1ySkPPxpEdn+CdIc9BVUEc0Tn4ju44c4AEBr3Og
YYS+kIB+0S+3mRQ3I0miWlP3RV66T7r2nx8ggT1RJzbsIdYU3prSqEJdiF6RknXo
qKg8pJpR6oHgxDslKsuSYoQCo04+M8PIEKeK72BZ3DF3rIiDNkvK1V5RvaNPTDis
i/xQQ7QMebomnvmo/kjT7E9frcN0VMSyo/bfbjZf3Yc5iQ8lXOQaUwpPs5fvufCi
7hODcApXg8lcZmfMcIjoUUQOkcFSPVqj0C4vxw8Y2tBJ36wRgKJz/O34twtde6pi
V4A1U4YBXFZp4NDC1T7rxhxb6T270iEVF29DAz8ylpwlVK7yrcq+eAjP48b29zhI
VgxXGbo1JHHl9FHEJ8YfagJaiIHvK8zY/jg2e8XyKTmIWM7ODDX5w/msiF//ETdj
5YBIR2uWZfJ+Nss4qRxFVhe0FiKtoMUOJGqFpEToMmJ5UthDpKHQYE0JbgFRUbIL
bJRy7YeQc95gru18tpIvCDiSUfCflXLN1ABCFAIIXR6pqS+4VZigndqD7PmbB2xD
5ot27eUe7MTeY3C4rxApIlf3Uzh/RW/YMvGtLUQxoofM7t1znp9vhZV4Rx1RjTJ9
cI7D2BVP4AHMFSt6/rzh2eOTjJLRQEJjbvTFbrgtScRSzt9Hs2OgeekemIfSJS9X
CvfNk6/E9c176mUEyWQUl1oxX2ZJm1dIbVTGD093KiChHqaZvaeoDU9MNiKdIvp2
epuw+7xhCYdB8pX1lEALtKJLwX6/0J2oUn0iuLawLyOUWpn7Z5novNtw0n0C7YQE
witYvpFFAvR0JnfUjdxqaoqo3W3eJKMXf7hsP6q+DD0AYfTpPCCzqiT1UKXpo9Ew
r0BLZ1IahvN6yr+RjvFvkctVnqPl1YI0ZN7HZM0hw+QGEEm9TgvYidYnSKpWSn+K
loFuoqhTKGccsM/MqfLkFPzuJ05vDoxCSKj2BhpouxtptNKNHc3GGv5nXS71a99e
fyinpFnKSmPCdDysGoNgLhuI7Aj+y+1wU03xg0RCFfxJODlgXRHbNMirP+07gi1t
PnfCnFs6Pf3xQkxxXeTE4Ioj5UED00ZmVqZrKa2h1TkNBCT+JY5Gy5S/5AjTsK1W
QhpaKJUhyYANHvkmp1E5lUSMPFsi+G0BkNpCN4GaAj5uVYZwv4jW2YX8YDQmMl8d
Tj7yzorla71LgoPCgm/N0ZgnZrk4sWM61XMO4FskK3XokG/rY2YWV6Tu+Fvcli2u
C2A8o0GT7L0Ve4pqzLSRXr7IJt9PAHwKPjxobC0pxQGhoXs3Ixe9Py+Hq5WFEAxR
wd1iHjTdlg0E5eB3FwFy6/8dBFxgvFExF+zB8Bqh2eU8vJo4uQEsLpxXuyYvvNGb
ocBZ0ytEHJ78hHxzVTN+7l4vZV1+OtwM9MI7ZA3cR/+lXESEdygEUpaGSDofw2fS
c/g6ytQqVXX8GT6jBKs72eCS+uC249eup8+y4np39F8Vob6ASGULTDaOS1I8/cOs
VL/JJWduPKs3EYLSm8PO9kDZWUsjTQjWBklnaeSUnszN9WZl72H7njnuktadpB28
ab8yHyVb28/hDzhEcNjG/olyFRKfODG8lIoFHuBuybNHztwpca6Gi24/jISl9bnP
pwsApH9NFbzt1X6DG9cY77cNvzCL1KjszI5O7sV/aP+KkO579RoER1VzUIj1orew
HrVtPhPb8VDd2b2LV2ZsVFNsgXDZDG403cfnHOrxIQgCz8/2kilZdy8oLFHummRI
1GGpOo8Pf7M38+1XKjp+S0ngFkfrf6AJh5YahOl+/38tZvlGI3jQps+uHM0viQ7V
KP2zQEmJ+dYXjq3cIsBiO27iX5NynUlA9ENCNEy51j2WGP2RC+1xctg5F9U2oskG
IwFpowm8wjb/rOWvf1JayKyJqH38X2hxJPcmt3leBgR3ynNjxSlJ+PVW3cSkv7ua
O57khM0zp1pAPsJM6U+dxhebnG6/tJiostlgCWmDjqWals0RLjCMevtK3T/gVygG
kzLe7RVH9SH88aTzRl6LLucvDrk4hT9WBmA7hlYRQVsQJcBXm1OkzBAK5xsuL0A8
SeRLkxxX4MjC02U/wuTmckl0VDhqeqGF9tcb61/TVOl3VHUtU+4xS1k3jXfsB2Yo
XHA3FkGHdovORLxrpxCYuQAhXQA0y7nfxWmm5MTCLOfNACLWJjIJvszWwdok/BLw
jtZnv4hDW7y1EyPxXsSmdJFdbs3qorJbJyBZufo+Q7oPS6ue+QBo8I75kaAPpotS
0SZm4OR1IVXnobi4uQzzKr73ftTcBD0tJBybwqbUMJP6PgtF+9vAYAWUM/dRS2Y1
8Z5v33TqnfYpTWtQbwdz2PhkQEDl7atBWyYpgylo9horo/OHOh7xfhpO9RO9+38h
9lKDVxysYaUI0HoMHHDs+iRIsPlNDRc5xTcoEGHW9M3VMGfwV7FRu7z37JmmcIdr
xi+j80PvjMwRzYTBkQPRUGh9IT68yr7Rxaq3ydLT179bSSpuckSVHW/t7rmi0e9H
IW+ghn+7+zvjcUbA/im+XoGLg6BSve50x3px0RUJG7tQRMekQvB/GY3iLAHOSVqn
EZUYPCNa1s0Pha+hplhahOIpIgy/PZGHItVdWetnKYbTlIvAfxPeu9df/CRqZeoA
YbXlRiAJvDihX2dCIfKJh7TLNctVz+ZisiPqzKbNY6961BpYuSvTYPWShgbmQfdl
EHNP7JkNYEoSwAbhoHyzDrno25nEdi7CoeApC5k20ToNJAt6o2JOz4f+x9qGdARL
UKa/+4df1Rgszdt137b0ZYfUPn3DpYkfnSTezFxIKF6r7GEJCO/uKzUdNKRvGtda
HTSO6aOcT1gCEo+K7Nw9Y5Nm6cc/EsJVWE/iUgPl+umI0QnT5hfdwicO+VZSoTQN
IP6/jS8bZan5pNDaUNyl2YPu3slOrpJpAnAgWGr2PtoLT/8aYamkniEGet6gAjM+
HK2oBbPu3n67OOjGGOJyR6XbK1G6cMIwvIKjl0f/N4UxNmuoLaNRP9HDhIxKG10w
3AezWkpB8iTsB3SjJsTfGWOcRPCUD/Tgqw17HDW8GRIq3xVA/Jvk9p4bha/wHjgu
/TvqU2KFlQFI3ThYtJ6/kjqTNojDVo2XtIuD3oadwOtUpUmS3rAIxJYI8svDpUme
XJ3DwBIwNVJdIzNeMWnm8fmT1WDJVRQVW7cGXMFWHdk+4VSWTyZbe697XrplyUNB
2qLpcD1M1Pay0JWiKg5BIJV4HR4SbzboGMHAQnjeLf89o5QM5DljGpZwmAd0NT1n
6ZVe4WPX+uu8i2OHC6qWs6lW2NfjZJN1cyJXxOUzYFy6Zvg/fL1kKUlb91LGXH/U
y2FcEP1BO0791+Yr0Ibuwvdc9XlIqeBLYjE2AFhu75T37uG6l4f8UC9DxUANeeMP
LCxZ0BWYFaTZ4cDlbIYFL/cs8K2xO9MmOYZ0qOpEvP3I5F6IOg2nJJThVWL43gMr
20JRyh7nvKiAGU7ZTWq/qHmh8Pp/Yn3elfJvlS6PdMxUnI990YcRc8iRw6iRKCDR
EVoodBeiigSqN6kEsN0uZdqVp8Rr8XZMnzB3zfXwCOlhfomOR2SCYnmXDXYEnKc5
PDYAyMYuhcWPp/B5acetBFPIhrikaUaqwt6U8sMYLJTyfzP4yRx2vPOYQd+Acw4+
6UJwoSUojHUcLltevzgQPjSZuXG67yHTxB/iq8hpvZKQT69SNtxmXLfHfb/cyiZn
uUCAJ2KmG68tCPNSbRmy7jFVYvyQ11WSUjeiJl/X0NZtAmFU7SkXTNEpzgcsGW2e
ZRujGNKG677Nxvcw8iMEw4VqiruRNZRSB6MA3Qe88PPO+ZqD9o+hjNkDK8cJCslI
zWA5g15tBL8bxt1d/uE1nqDmP7Mr1kUExSAExirV/qsOdYi2TvDiG6F1N63palNz
KnHLE5f6xXxmTG0xjZrHWPUGBZfKNkkXzSx7K02xAch8vHyqQUEf5RbYIQ3nsMgP
Dib0B23DZDQpgT9guNuuVOOXHUA6bI0I9get7IDNJ8/fQVZSaPghhNv8LxHmWwta
mNAtNGBWjR9AsnSVBdxXcjroebeGVAhRoy832w2S3tjTX9kSB+EYSHq2PFUOuYdp
ItqneQIZY3+XuGZpVKrYCWB96Gj4lc/Y9gtM/q5B5SbpsNb7ysS2nOwK2ekiFr2Z
ZPgFoD2DLNI20xWTFwbpnVaj7oGpuqAMOyVV3Z7Op73DIkuWHRKpDvWehJOUHmHi
LwjJvYbsNtjt5cySs7KQuWmCLKL1xFZa66IeU5a1IGr7Mz0wdqk1Chx7yiOJRR77
Wh2NXd3VEa8dwY7s3EMwWF4ZweivjBz/H6NjjdRqWwqzzBgzZBYh0l54iVkL86O2
ZDb5Qc0dDJwpzbTIvOShFTloIw1JRPgQsZvRnqQN/jH/pizooJP4YPo6Oc7Zzgcv
OJ8FMpQNfUWz3dspLaIFffy6Pz0nCoNA9bcN1wUPJvjSRqdm138hGlX7Wz89VnZM
dzoLs3lLKrisiCsf+aeoLxEaz92LmoAoE99vWVt58IyolQDP2vNj3cvw+9dzXc00
zee/QMkvXe4NculOieXeM5BkNbnxTJKSisHK88h8QIwOTGFLgrxKUK6lcVzrTB9K
ilqfgImx7O21x9kOvbRtZk1B7r9pGS4Xd4J30Dgz7U6iKIKWCkyP4O2z2/TjLksm
rEazjz4Bt8I06DZfFWmQPPcjUNxmpG263oSEcTtGtnCCzSAKWoheDYQfQ3//O17x
b0oz1mKI1llyJ/ZlNtPi2fg4PoVIyAZ1hDKxsWSfiIQD4bYWAJkpbb69QlxyHsPC
2qbgF9gYkDrVQrf2iSa7kJiNbgP7NoReZiH/+WGCEQUMsvFU21O3/pU41jqDaLet
mUUjq7xp1Iah90IgdFzqraXHpilnR5In2AKZxzJF3oURf7izNDq76i4fENkM1yc/
RC1cS6BpT1HWyv1L4//nu5j52xt5gBoXQO3HPq3YJwKbL/WoJOtWzW5fjAs9K/RI
C63RgVxYhaJh2SKo9nBtyJuFlEwAi/0a1vVhCtuXApKTxMER6Mx0VPooXQUnOcYZ
4+OUacZZ+ObWMkqJAO0a1PeN0kp6RH8CjqP2BQLNyKsKoCf6fUL/ccqj3vKV0a/d
05gOjIAMQ5KIQR6hp2ofcBe2xfRhv8KClGTR9NP9cnUoI7kiniTL5t+Pqm6+6KGo
5aTzWWM8FoX2YI/gyDFGh8DkpJeLZ4IJyRhcaIZdTnZHMVCurSPgvsTMun4dfp6C
eiiMA7SnutloBvQLduko9KIlKShcNHxcz6mvhhB+/ZVOJdzEOs7AJ8OPYsdQojq/
7Bki3ShDo5wqJH3613p5ofNgRuZDcu+sFsjKWi4w6tA7bXfKSUSaZAzdnk26ktK/
KaIuShfznamke5PB1hUyCdhbABHCT9xGjermm4Q5KpldzZffXO5ssp4VtmggfqJE
I25NdfnhIUeOGYrjFffsyua1UeRL/8mJOjDF2rPUneFsleANogR8zhc17G1XQBO3
8j8q72qPNEw2KclT9MippvCKvHeUay8cbdhHs+puq7FAuNMvWpVY1mHogbO8L/cr
/W0a5Ew87QB/CsVlBBbGiySwoCsolkufWUt9wcP0IyRxdmOw/29FImkuqSNl+krm
YmqRiK2mRYEgbe9y1RLoVibd76rqndgf9jAwBTQtwo2cWQK6FdOksXKTzgebMDL5
aj2g1+9sQWPFjLBnMm2DMGlPGcYSX0v05zRIq6RoSUN3XhmqRfBbJISz05Opm/Bc
nLnVkWSJvU3hwqDJcro92PjtO/ko+Hg6I4maYWVq8iaaLutbku28f4zSaKM8f3y1
X/+0siMdjbMRGnQB4L/iTNAJN1/xAvitemGp18vKLgkaUNvmqrr77UHzgXKOZ5Ms
9QgknhlNqKItXdrmZXWwZ2eCcKgRHTSzPO0XHHgkP+BluwkTqh5mwnDN6OMGBMxy
UPd3AC+rM5APGeE1PtpNa5aR7UgVgsPoxu0+hjguY9nqL/ojCSkcicZtSanqmyJG
ptCw+Kl300fYTRLX2yUHWdYsva/gKIsGlNh0LcoGjpTGxqosYaxSF0P5zpaPO+Ds
R5aW17wiq5Vk7Xt3gzWUnh+nTn56AYHP5MPRxrjIRr5nkhFZjPDlh0MmYzK7XA+A
NgZDlzXEpwzgTkt6ByP+cXQa6Axq+yfnJxJY6oWRu3W5WLfJ43UnLeUt48lJduhb
AJwPoGZJOzcTWt4ksWgYrnPQx9e31B2ikomh60ISfgN3b2eOnGPsy7/pBKJa/Bbi
+LnryPJrfExaVWKfmxs0FyO503HXk5Vg+2Mg0K6LZupCEZcSu5xGfZSW//CijTkZ
oyEmYMkq3jgXh1FWNDcJ+1ter7V1g8lp32VQ6afUp+Lj/A1XlU/g3/ZIrzhvVPXx
OVxCYukjLuN5DyyFdrbb0bUVuJ++RXsqjPO6pZHpLQYX7Lbenz5ynU/rkyGrZ9Rv
ZqfghwavBmjhJnRGT1v/uLPeEpfCjt5nCHMYjpA1Nvq43Glui9k7h9Ji8NOosMf4
WP+0OWgeW71FA5BPPt/v5oZBnA5fWLo7yLFcCDQFkDUenMPoh1K17JO811U2de5W
je2E9gZyS8MPr/gCK+TGh/pADJJVxMZ4xJKerUR37ARDAL5McOLxdzGpgzx/41JE
KzZbrV8xG6/LeBeGkxP7cAjs5U5UFUpZxXjTCHR3TV0XSjbgg3H0oijSBpiWrEdN
KDNQ4vHKiInm3FPp+t52T5NV/Foovq7xeNZFN3WRWS7qGSUawY/kMUkokJv4HenL
hqh7ZvBQOKiNOGXHo7s0/Z+YtCfFm4EYJLtxkbcWHXABMzQyPF4Hh2MWtL52FIT5
JgivO6XuWRxJhbYe4+DVqpzaT7u9dSlzAKlhLhNos4+i6o4Zed3xE6Bg/DsLmZjz
3CSfCsFd06y/tMDThR2+GVEZBUmSod+u4v2X/vDWm6oG/MBLQheBsFpiJnUgHmbW
GQz300KcQOpDKhSac8eDyZaFzYv9CbiAsVSxeVq1i0KvI1VnvaecDwTww2+TLQsT
sps9UFVOrX3zwtjpEFnufqCalaMK/+siwut69aMv/+XbfwUMIzBCyF73mkIPoDlw
MJy3ndDlKCAvLtF3Pu93llBrkNsvv/1LkB60N0ITWE3UWgCijwLnfeXPjg0GakUI
K2HQyVUm/V0L/ZIupOXDTL/QshWE0i4I9eZAjHh9n0uP+eYSv8U+RdOOgR2Ho6wl
s8AmACaYP1w102FuOq+HaNqh6cu2wr4sLAOh5ZXjEPmZUqmPAbSd1aumeau0KQ7G
BJuZgxtXJwsTKohfj+/PRb39U7/zQuMCXcXP6lzWPHIdeP1kr658Zl3UJQX/KERh
P/n23OPAVXXWNd0xjKu93izdbDzetpsS7EPxhnilbGnMay0nOoqleS+P+EG54Tjd
ZzYNkpDxqU6dRuZwl0VNM07vTvzZCModWmTpQtxm1s6TLLTxLhRdUsVQ6+TJTvPC
/aEokKhEAW9+Y6XWcIVeHH6dKNzRUWSUwWvQ0OIdkTI3zxpFuBu7iLD2B9ktLqC+
e7AjzgCF8wCjck0vX0TBtwAfWdfDneGkSoYhPw/f9hJMpR3yAHkgnDUGJDh7I/YV
S/ymctRgr0RR0RH0Cg7QdxTwraCiyQTBViSWg8/rKl5JisHx4amAA9UXEJbqACZr
cG/IAS2ZcgBZ607G/8vRp9h12Nyet+eVzumgPzQb0IU2ha4+9WQlt4+PC2xNCcn+
Em/N63yDd2k9lycIzeoHlXIKbsNx4uy4NzPuNUYS6Ke3iIygvZUYJp95nMHIfALc
H5JyOaDYu6jE9WifZ25o3KR+w8lZrYkPbpyyT4F44lihbi9MybyDo8uPkYzfZNKo
gLF498Um0NN6YQocSsrQ4zaLqtI4Oi6Zo9SetQe5zKCefTVEPRbkGu5xHbLgChY8
QeWrnCQwL09PTc2HlXWWTuBeQXtDh1RomSXnuHIW3R5UxbkELzdu42bOmviv6Miw
lxf2QknaNrcay2p3u1T6KJ7LGyeW3r9SkpmBUEV/WeghzpOUdgj/s4Vvc4C2Rejs
gqtjXIJjf17ssbAzmZTjVLnY8ANEt8J/wRwAYdudke21UOQxUk0G0xTugeD0bknk
xk/7LAzePL89dG4jLT3bRdFX4O+dkBJ2VAVZfiEfkOdVxHNCyO4IAXfuwT6GVI0F
NxS3mpkDuBww+/VliVpEMTi3fPwvBRGSrSsp/7JSLC05iXjtZzwnGtxMc7xv7U7h
/ByJwRQWeSkt03VZtF5VCXU2k/O5wYiPw0LpqahPAMtC2sfGtIP5igFfR+juG6Zj
m96Ue0bIjOvRrISR+iZtohsyGe6YME90Jj8+koOys9mX4YDvn0Auz0j7kLHqUD1E
cNczxao/GxT+BAVJrtqHcCASGe/FN16MFdI7spbmAI/HE76O+rpG2P05IW6D+STj
/TCi9kWuPrjIX8k4uTDX8RqFayqX5FMwTurgY4UrMIJOqU2gJl3K3PM7xAQuOXnL
xjD/InBmcYQvVJ5OHjdgFuLUFWdlHCCQa59B0AaFBospIJwCVUzWvz8MLBAobOkf
DRx57vnoi+IwzXiwDXmtJN98wD9JowuF/OXf0ea295ZC0x/ze1W1K7NWr3HfIOk1
dDHqFqfMfIfUW02gLnRdq26Xd0LGhwe0LjNhZU3N4NLjbo9kWPEr60jj2Pph+7Nu
RlGkL/k25sRN8ZzhAd0rsJlnfIh1Gkbj7wLPMQOiokjxiqzH9wEgHguh5VGeJnKu
NtpnX8Ay54/otLRfiAnW38oeX1Gy5fmG0sAZb57+pCxt/UwaDmoUYXR0RmVFvQ6f
KcACtOcLX6k4kwhffz9K3RE/cK/16YHeCWXQ1p6CBtYWeqPGPqtk3VP/GpTdEcBw
rPk52fXV7/H647tVj+2HuHeEKsh+7N/+bFovuRAx6iruLT2D5Qz500XTFS3KO18S
e8n2Nmdl5Tz1NUPiyYkx3OQFoWpw2aWYP7M5jVNSrWcWjXK3uxrmYrwOJa9ZMCKm
uSZ6AuiRdNwkRQtAp6OBV4wmyV/ERRI//jPze7OL7nPhvyE3WRcB3qFHv+0rwAG2
I8yH4AuxRAW2A+Ak5h/4ypoo2LAqLJIQc4q8i2uHbG21XNYrtoAtyczeXvEUM77V
UtHlwDBjuBzg6iNGHm8CDxT0UCoc8quLoS6jCQV3qjuy2QFjKCU1CWHtlokCpEtI
pRIIG0F716h5xmWyL9AKBVfoU5C/qPX4hpcsfwVNVsR0xregCtp4Vd5ldKdwGnMX
yusS/ed/3Tl0fkoEqlnrrzxZ9uBYLwnw0MC1rODblJ22TJ7B4VBmcnt9giU9OmK8
lPJfQEnHVltwRgG3qQidfKNT5RpbjlJvmXyqwRUIGLduO00a/EdGMbHKygsSybR4
/ZwK2e9rxKCkqgPT2E9XTrxrC19zOhbuq1n9MSJ8X83B2XE82HJVSYQ8ojy8/U8a
2gT0oItwMvCv8mbGwLokee3JTsR0ebsiKrAqNrmlrpKQ3kOs5HJlU1J1AP0mVhIg
TqmQCNnUeQrgikk6Lw1tvW4BP5mdYUholXtdUBLGj3c58AjL3R2KlTquimkcPhQi
BAQHwbJiaEdNcEudzXsMda0ZqWHWatYHxUGw2SwjTJWYgVTLawhrPkB2DtUnTS9L
nEvu4/sBX7WhidPU2Dolcvh5ZjdlBbVaU1hgJ8OI4mZfuXvBit5DbPB/U2hu7bBw
tayctmc8V6GXxQI2Ht4WTBoAUqtYELwJ03xly2KcwgmYtKevWerUqsvCt3JKq18z
uc9SXUn5azJ+5HJiNOEuzZo4DYJkZGAxERXDafU9mH2Pyi3K36Scl+MtEU6Z1wBf
vRP/aD2QmKA5iAUDVjzkjq15N+p5Hs23ruZNY3LKKq9Xlbvy+7DaHR03YSUFCdKS
zIxle9FaTawo6dsr6iY14MGcvrSh8ihkTBohkm61l2Eze3mfnUZDHOJl5iYq3brx
R8fbpndo7CrsT8QixeMtNqFxtnUA9T4rqL35E763giSNa3IDCnLnn2uKcBbDEiNG
UQ56IzzlhoTIuYmZMONBGqvbUYkHyFcEZWeOK7DuUYtvLA/MjbH5l0XxRpxWQVA5
yhtbwHKBphd9xwSu/47e2qURlsgmiTGgEa/Hlny/Wwk9iiwhwvB42XvaaLZZxJU7
gDy0cNpR/V/BgBppLBOAesdjPbNVdcWb0dkIWPeS4f3C/p+TErUVvjUZYifesTZg
W7r8P1c1GU9YTAy3Nfct1waBv9hZlhTXiSnmt8aEOT9eQHXbbB0gAkueiDtW159I
AR7FHc8pbBjqmZd+vPLJM2VUJoW/FfEREeb2pazGeP+1SwJH+dKB4ewuCan1cZlI
DFMWx7VF+X62yL1cUYVRHDV4kkGnPTcy44LOVIKUjlJkCiqDxub0Vn8567+LWEFl
ccPgTOGPqmje+WPzpsatdPhuaTWOX3SRAvV70xlsVi60WTKwlUD/SaXD1LTFMyQ0
LgbajrHHT/0XANqwe7ZPxCaKZMXzzi20vLzCIVkbwaM4+WOuCjh4X0IHjcaPLNM7
9m+7vvI6o5U4Dtn7iBuuaAnFQ34IB1v5jqNhVDR0kWIDym1UZZWb3YslOYPu4/Hf
FUuE33mW+x7m9r7tF8/hSHVuFlhOJ5vfasYbCH2ll6ByphAz/NaNRwMMhI/4/A4C
k1wW2pUYNyqUKy+r/aNEryTB6cCDhOEexOF4tRheDUZ59Y66R29dfb5fZtAQXWwN
BW8q6GTgI4/bXEPxeZts8Zr4VaQgX3fQf27PG6XggIysf0NzW7j9FxcSr2KqKZkw
xOs6b8qMNf5Rt7x4taor0gsFsWkVlaCOmMXbzbUjnwb+N8SNKdTlr94Sauzk9jiJ
5nDDjtS7Z4Rp7Dhe06vhcOE+Cm3ORreKO3NDQjIr3ycUPE8sFpAb09IPJOmPSuin
vcNqEl7hzj9ASRyetpuO0xlLz/H0Jr7o2GvZs/WSsfyK39Y+aoznNtdItYi+AA5W
/KryNRETwz1vJrKPlcQBh1HF2voAk+P3J+6XHP070ikXchGMP+5KpYlz6sG1+UiK
qJJEIi7WjdwL9Lk31gcCK90IGc2hybsyjq2NfhbbbwOMQb3UvVHTYGsO4Md1oTCJ
gVf65UfI0dVTPL3/v7OCCauofv9okvCOfrssr3JM47WanWyvHC3usMd2GYHTnujb
TsDyUnKEoaNFx0PEIEsbBjS0PpGTLvdhPlA9Wze2ctVaVpaJYNfxkYkfjs8Nt3yX
wus9AtmWVeIqlNsk9RkXR9FzI1u5Izlp84KW4rh0NT2fxEaQouqMqky/5pCEVkie
ZcayZwQFALPctFuTbsCckmgvTgr2t+hHzUXINVifqjO8jdini/wru+qv2o9jzvwg
VGML0CCU7pdHsrxw7/QCQ3020DKZcnRNXb9E6mFqgMhfHXOLZJYJBq2BJInTTTzZ
c2+oI1g1e/RWFkRaLECRkgraOqIIPw3rPBhss1GQ7QvuV4QPihSxf1vAo6MkgUI1
IXeL210JNxfHMU7yZolUkaXfa05NQMyLCWHkTr2i6VZKZIg8C1Vur89VSPFkAOFD
+mjdGIEd15PqlN0cKZUWXFxekAXGPG9Srd+2ERTn2O/G0fopO9BwtwTfYNPVkxtp
DauMDbzKPKw+JvlOGMbdGkktp9Rs2nvHBUFQ9MZ5STelHgK4oap0PKMgELQ9f3os
dSU8fryCpJDhrgbUoGPR40rqxHUxh7TlGG3rzjsZp1UopmlaA5lKJrtyV8LxRVF1
Vgvqb6qkfz0Ijd+r1bI4UVmt3rc44dktta8LQrefDfhFJBE02NmZ81SyGSn8ON0U
cZL0mHx0GD8+9w/pzyKSzyAP+9AqkUcPEIVEM9S1sLQTlylPyK58H+r9mW0xA1N+
jmCAfChmyiDAdwpzBY/sw/aKYRw6Oe89uavKEXa89ZsYYMtvgN6OCMigCkrrH2jV
C0XGAc94nkART6shSZPEp2JMgMh6Knky5AKNoNMlcXD6vqpy2wNbw3c5UjSuuPT1
Cjnou83TMs2h45X/Xv72DMHYJocpmAvnU+tBfrsw1MVY0o6dAwOpHGcX9WC8rdBQ
XdbU/GHqJYVQoPc6nIYoYtL5jEr6pSmbRZR/BpW+Jm6y480kQ9iewN5sJnVk8+sT
UpX7c5yHxE+o0QypnQhG8156T0yVXMwybOigGpwBKm1S4iqCdPzRV65Rv9QqcGQZ
u6FCFt2XsdemlB3RHABVL99AQ8n8tMZRuiFxbYhsHSSF9jxbFvCylIj+qzGBPKqm
2nRJtwUQ3sOlwfi/gzsgByHgF+f2nEo6ndme9rgxfC8pwuBZ+Q+rcyCf/FZfeBcE
AzHAp070OqtArX8Jlu/3Mwig3Y6R9ViEL6GhOQnTnc1zssABxCHafyjovMXphrse
G5G8dywGoEDRv0FLR1N6CdveKVdNWog5Ls8MKaTykHghwbY0PQJYq2B7Kq9MDpm1
PWq71RK/FqA4pJXpJFBB3PqUOmp6MC6zddOFmRG5S/r2BZgI50F0b+OcqCdY4Kd8
5fa45rht6Wkzq8lbM55fWWN5LOTmrClaxUvsUv1R99WadD0ut5Zcm9S/i2OViVAx
DjEujzbTLZ7ugWw6WxFRErxPVPWL++87auPn5E9odw4apT9fS3IxBWc/SkhRrA6k
0IlNqCHv9YW9EIztG5ibnWd7oyQT5/8U0r89aHojYwrl3waVePvjDcJmGpWDCrs+
ew4RZc+EcncclHP8g812rgerKPVBZaYH8mOB1oml1GoNdBN0qb057AX4o9fELWRr
Q3OQnyRbont0iT9z7zx33TEC81uwgm3qSj0WQWZkTf62j90fFGfZaTClo85BSCbK
0S1yBwacX5QllWO6EiAacko87TF78gAjv5GNNHqE/rne57RUqBUypT1LP+sfwGfZ
ary1qj5CYE3k3olWQ0T+a/ecJodj+P6QaktUYSIM3k92Lvd1L9522dFlckETAhh6
iKMVGksgzs9HrhLql6v6GZUTaEy9zwTC//soNWUDr5c956IwvCvH9x6C4hI+ZhNV
2xeH2PFetRr8v3/BBPpEsirgVN9PAOIXq3fGKgspBGNsHQhsx32MgGGCn5RmdH6j
zm2VZbY4l/GvcrS++pgMAdQskVEPHC+BSxSqdJbbjbBvoJbHaQdnf98uz0wsZ1mW
BjUSKIg/qqqULY06Rixx0MiTB6ONqFvfiE4W7gDYZK+aD/aU65jyEefiU1YHkjex
iJqGvNkJlf5GjT8HwunI6sYgf0qYKGd6Cjt81v7RXojXG176AAfs+QTARLKLfxJC
FEY35VKxNIa1ix7Sg+s630tzuwQVfwFejTMSw65eFutQg7DftgYJXazGr7bH7J8S
hN9dbchrNu0dl2HCOGwqLYRr7adJuKsJwq74xLdbxUfZQay/oEpuyfIf2WSrDMFI
9XY4w/QcQ/FcCliEyDLh4kI3h1TELe3Oa/29Y8kvWd9qs2M2AP5Q8OeoiOpmJj+J
+jttwXesed975R6DsJoTt3BlaDHYKHjG2qlLxn1TTJswKQ9ukp4AtRqTwd0tkIfn
l57RhAJXkDPnWeTDLhH32Y7C/QFYpQ2BXvYZZOjXGc75j85Yg4WjpdjpM1on8CSm
R/akSAMsHyVafdC1XJcJRV1b5eQPlJyR8RpXVp2pgcfUdUNWEB/TWvcrL1vRNVo0
7XhwZxdzVm0sv5Y7oRzEeOiJIA2POlkVsHLYjKC92AUEMmC7KrGFN0gi/uvmPNAI
/yLGuqgBVRtlDy9Th8X2GDWzavJfDuPHnRav5NzlRe+sc0LUlF3VHGOH84PTTHBM
AavQ4P2hgDme+fNWrE3e1c/gWbBTc7+6kIs6gpUdLQZhsGjZDzerju0V56tgDR3M
WRE0qgv4YWf4W7OlJKlepXpuNuYY3MXEXCcMJao5DjXk1R3CGc7knfHyHJDWGdJh
4o9Njx3EMTv3STbeDa3z6kt09iT8fngKG1aJD0c+CMwvBeffywgYsxrlUIZc2NIg
BmZd5G3ViNzmaT4tu8UomXDroCZ0zFqIUTjUqw/GBAxi9Fi6YUhYvEU6gDe9Bvwy
FAW1qdg8SGNQpcM90NwkWeTKabYASzfmWKgTqzYZWaIUr5qMcyPfVtULC5LQGh4w
8r3OB0szkwST2XZHGSQAWY33wcshhD9ir8cJWyzuBIdgKMfU0IxhZEvtkLw3bhDr
MU2vzh8Xa3LS37R8jJOXuNTStAzMBPT7trGAx7H1jVJ7D+J6PAl4XhgQvC3YBH8r
2A0YEWGCJljlqdrgKo7YUlKXMlNBYNhuy8kCCxKNA78Rux3gof4ZqS9GBDhYAZre
VSnA3/CpxLE62GlE56PZCizDAx7dQBYMuf8uIQ4OXj3gj9vnj6EIgxm5LmBbUjC6
Jf/4OCdNJHzuATV1cuI/9f8VQe9Pktz4QHQBiGby/52CFnXRU8kNKPFkWGHlB4Or
gQWerI3WYJUnymmu9cYZZ8E5JJSN2+PgU1LOkXVqAxBciukurvzpKmdq7tlqxir6
bya3AAUc5drfcgAtag1jN9tOMkaRq48Wo/2SWdMESxffZFX67Rj6BYredFVodwGL
LGu0tJy/aGv2Ug5sCwXAD6o8m5kLj7wxdyE4ln5mBbhhbepJ8XLZ213JwJ7BQA0q
KPOwWFsVJMceHDwHdXq7PPmkw5YzSaiaNgkqxXClH8AyzybfpCxHGSKpAz77WwIJ
i0LdFDVsGY/7NkttBVc75X1+iRKb4dTMe5eR37xCN1FzHOzk/hJwt5W8y+PKHqiL
WL029VaS1z77UDYtzQKPL6FradPa6DkMqr3s1DrwN7ipGi1fymqFSTlQNnkCh4zK
687Hln52va5gUV6v880+ccLdPxNwKzRNfgtx/HQptdSYGcoUP+u5hcg9KrNvZJG7
kUhRfIpH4ROzD9P6pxsRDgl3Ycf9Hea1diQSpg0CYxPfRosEPTxVWxQ0onbqXPAt
vI2HFHTosNPtIwgBiQw0rnwDZfQl1FFiVRsFHxWsDi8IvF9xdHmUqOHO8rGYVp9D
FxCCTLhojRGs09fyyld+ywgBmylQL9iAz9yt1+ADpeVgCQc5btmWME646hy0a2dB
9vJIKSyzfWhwPF3+s2Dze9m+PuP9T1u50GbkHVRJBhG3Dy1i6dWAO+a5C5YBhQaF
bTs4hqL/FbyAoWSSGMocoAC+yn85kiAVbkGnCymmo6ZWbg9JuSRhfjdJoqPtxTDj
BGxjoKfCjKcYNoqr3OTwg+HmF5ofXV8XsCAJzyCBpkm4uAV2lG1JAzPmsgBXEU9T
scjXeeu///aprDazuhjlkxC8x1PJvtSrpxXuhceYe6vbNEWh1nWa+7K2oGUUNCyJ
HEkHOBPK6duW/atx2qep1FZkPVr1JTefLz7OvuAsjGoz7GVirB6KfsMxV9dKVGux
UFSETlP3e/fvlj40FLs0Ld8sfCjb2A9GPBn64pLjngmtS8cRHSCkFF0oi1X80DLd
EsL3c6qQNhvgYwJA6OqXrdBDrTYyIgY2KYmZrJ6+LeI/08vKL/WGeYIAQZPsWnMx
1hO+nM+eNQMKXsaUQEEIajs+h4KSxjGSwp4tZEtebpy7Y/XmzzOcwLurd3/zR3UP
hcaGhOg5BchJZdMCYRAnTfdLm40moYBOhEkwnmfFxlwT7gBIGYlyWWk/ECtzA1Yp
i+DVeFgfa6sQDlZmcSKZCtop+OSr+6aY3k9Buc9hwcRfM0RLIl/ibqSOx5791i6N
dPnCXWg+Wa3y/uAqkNVLA0lSfqaueJ20kXIxIVLz8tDtbcttLG/MAWq17rPsvQM8
Dwr9QldpHG2MPkcCPqpc11GIMkjnqnGQkAgiI7dHZVS1oc0CsHUQmW6/MeSxe5+X
zZp2lX3EVHBhiBOi6XQMvXl1ltY9BcQLw/0pmHE6aRbemxyVXC+SVyou9xa/upLq
9ilHeabiU088LHxXmR7D+OrtXNY3Yl7R+xNvgUG5u4U72i74y7bKv6Q6bRHGzBIu
iqDfv8jyzjIg9Ks3bAsmKFtkKECjr1Y6nOzDIcTEnvcQr/Old62720j/DG2GOH0H
UKJf1m945vp6/G/9K7qe4UK72gCF4ny1DpJYnhjlsW3Tmauv+Tccc4XNAedjk9j3
ZADm8SDgVTf5YhNjUyOiYhXBE/wPHPq/IscOOmWNJt7O4U21D0D+Gkhrv03pKeQX
lNwxwcVIybjNtKuKNDJSMwAhcDxgktXjFn+WtRuaKvZPc6O2JgBvDR3lvPR33+PT
Kk8UFy4Y7G/xBconcLiRHw0bX/U9TJ0yvYqmGdJ2uEN0ehM5DgiRoREUPHZid88J
qlH+fv+vdjIpQfITGui2UMJeW43dOBFvB1bsvZKtfMjSXt2jtNVeICYu5EcwLu7a
0ktk2Cpu3Shb01ezB6LgX+pAPKPsCQmbD2lXBLlJKXAw/Ln9C+5t94LZyeoCl+UO
9SOwUNqaOumuPixayetPPNYiRgqDrpIOcN/LS5weVRmNKpGmw5xYwAQy4yLG0Vpl
RR+ArIwuF71MEx9I0x6yUpCKNOY6ZyyQAcrXurPyhalQg8lnvs0SV3S0y6P0pINy
LXk3MyVFY/1YZrl/hwTlSLDAxcPvogPFwfj3wjeLoOWu/F6peZysFHny4HzDNMjL
vgdOc5ATq5R514inFK4iN2fHUkuUURldRh27UfcMGmcFGWADyeKo6vHr7T1Lc0GL
8QogR/ynIp56Sf0aqmby9UFg+idDbGJOu8rXUaj65REH0hLXAFk0EgHiwFXQvtIu
PEMXL7UchP8N3xcQ8c5GTHL/R+y8EqpPFwAcu/cdkNUn05dZtOBy6te27Zap0mt5
Qlms4eHRnICnXlQ7+ZeMg2cWlWStR84cNxARMQCSqCxFunoxCDWJVnHYbhQRtgdY
IAxLfqiZos6GDeSVoNsuYDrdyibxCTOa5AG4NZ8jzzIVDhicsLFF1dCBqsDjT5xu
dGJFOVFa7Fk2DsbCQQxhO3lrs6AF0khZWPaTAqTG8r60CYk+zRI6R6R4ovWdp2cq
tQ1b/Iwq9tQpLiujitLfQ4jGjJEIZkoCWCyxSThgxprNkvHLUYxir7HZtyA7/QPR
Qpqg+iqPqZ/s4gaXBpF8AXd6zR/rgj9LS9ZjmDw5of/Zq9FS/kWzSq2y9Zcgsvsc
gnbBQDs6P5qvk3CI4/ouFjEKvkkzYFMSTduxHBxVShVdTrxFRNUTGqy/l52Mo8w+
03Oly0wCw12tPNQpTzTSVEjI0ofaAp5xXOnj/ijw4DqjuxqitYmKkGxLBgOT5LSw
AZF6Oxw/q0XmSyaJc6AagwXAV1yG2qbcyv52IlhGzCr8/CUB2vwqlV8kt1NwBO3V
wP3Wa5hy4/XU9m9LGC1EevW70RDh5ug5iGh0dZ0rtvVzoAqAO/2DAHNKUx98SfRO
cpeexKxrlGqvd9ta0kN3fqvpiEpDBNY828tRjZS7/yKthmE/wjD615IM19GYPrt9
Z3KTgtyj0+8I4z4D8O9ooK9QVb/9iTgbyrqhqOmA0YpGW/1SZb5Pcu8R74BcUWHz
xGILYkGKeDpp5b8zmf1+TYmPWBHSndyus0NzUamyEhWPNGxzbFfrJVj9Qfyp4Bas
rgpN+cPfDULqSi5OHdHzby6x4Txz5GpVDK9xJGyp1DReJic54aUk5yJ/RFKqzneU
mCIZipWGwh1ZRgB6UqV0TEJopxNRUc+9dWrujzhMKUg2fP3XCiHtD6oyEn3JQomG
dqzTG4tNFIyTyiqFiCgDo+/Zz+8vl18OT68dodXcOwVCpF8mmjpluJa2ifRaNzja
TOaXlHO/4k9Zqa40eeFaa9qEiu11/BhLGLTfyWVyW14mJTQQH6XtSfoMj5a/+sc8
CCfSZY36aW1x4SutW6kYnLQpIHRT2BgI+Fv1pwJUCpIYk7fkPAeD8fSPsKsIYeeL
7hE8ASjt9uV6l5y5sAgtymbQB2J6HrX5rHk8KFFDMqjak3b8Mi3lcHBs6C+gkWTo
ufKWm1hNwGhi9hoFfaW6GP23n+WhFFVYNdTdeLIvAQzAPldadLdZBNmrfAAWhYB6
Ew3h++4XW2i6g4uwaNnEr4SSHxCNiUyZh7jxyOebZIWpNIlgCr5kyHQMafuokERB
VOhPOShpNhwFd1ysy81Y0AwM+sFdv4ux3YCGDR7uZ8cPvN6yJpptQKacauCKF9nq
i5CJtZPRUcQOhLxlZoEyIpmOxHnQ9dLU2c7CnQUXLdHpC/SIRUDYqXaRIdOYsixU
H6LlATakcD6wLJy73nj6uCE/xSYEl37Ve1QnOT2Xow1vQTXQ83ph85DJdSjUwmha
cwuEHhJLGQ4/+8zlelAFtq13JBW9nkC+cUeWB6mST2V0fY2IhETm7nYTqDMfSeXG
hmpaG+O7fh9d48NkyT3OCFjmUJrS7V/9s3vXw3NW0lEAEUj9mDvJdzAA/cxC/6EZ
LD7qabWymiwBzemWl7jWNT1mGFPY/FC24IUwExwjRwr5zOWyJM59I1bmwF7Bm986
IiRuWhYqq4XjJkQr2iKQh2Fd7jjya1pDrUTwyoDmFhjzeosg4YOFge7PFSp0KfHe
EKZj2ASjdYyhmPc7GkYkihLew925Ij0HoXooEQQ1/dHZB7Su0eKOtcl3UopEHfyo
sFFr8H6HAzTht5NcOUWvBTX0tNCJ5HwX4B99hmuTgeAxqek+gjm+kRiFASjTsiBv
YhSPynH62pB+CGdaQnL6kFhsGXSO7i6r/b39tJmn8ACUpiAtmhRvakTeejNv1LGP
R29hMO9xMMUd4+niWaeitsO+r3+4ssJQ5GeluRF3aNUmETXY4Yz/Zw4rluMJGwif
K40uerdX4TWwtnMTJs/1JbzpVo+q7/AHqQUBpH9jrOfgIZ1+eOEkHA/OrJBQx0O7
4jc6ce3mKjLlmH3oQ1gqq/GF6604Iqa9JgF1PlppigbikxFqoogoe77AjKYEEXrO
4fm0bRpFeSmim/wM2xoxr6XdHQax/RcvrKSBDyQe3FVQNUxv1ymE1esaMQy6Z/Zj
Q4ZMSBDXXHdoPaNPmmUSWst5tFGHHu+uDAG98jQagF5E1r2RGn4BFZjHR9tXwyPU
Bzz9MCm+OVAFBfwU3aEPjDwtKH9Qq83gS+qZYR4wlyzSt1ZuoQmwdUaMmeghSQ5a
bE7SNHWf2Dpi7Ls44ZAgAhZKOBUcsrgmFAju1sKuHPjn1VBsCaT6UdeYslyjrqXM
N+wdY1IXEDMTgYcAA1cOaboJlSv+DiRFEuxNSfjeesD17u7e9DTETM6XZfopoFPJ
7Bjlam03nallqMJaoblWpmKTgcbQnQpaIyyB9IfcJ0qnjPgKCfR4WYBCFyuMY5VK
IGQiAXUd9OqfWUMVRuXbPmiUX064OYRmaw7ndABvr0ZKGCDbYuB71MW8wBaF2GEw
LbsBxBflmUwfLtGQvbnKRBitAC8R8C85zHaJjGWRYaXs/qdhXpfETgQWzmQ0+pGz
NZyVj/d1/1Qaorb8mZhKY/TqIvju2IsmGsok4+iWsCGze4fLeuw76yzSTb/XDZ4s
Sbn/qYYnZJ/WrLcgfFBVtWg2dnQ+axqVpncaDgDZFj/6U0r28uLWFVZxMzAdgjJx
dhb+bdksNj5Mj4bDp3+dJJLP0AmgFfJulEnEdMPA9cBvyaE2BlmKzFcxDJZr6UaG
54Bad91vqf2fD7k1eVTup9ZGKmYfiKxmNONRB7UmiDcpLwejGUgOvA+ICTZ+lD07
AAfIVHkSwaDZ9UQxNrky4eVXWrpqOyyqD6G0YCMhSEtcf6CnnzqlLXo+u9fdrkaX
8wyYIpuJ9v8xga7dSxMS4hfexNuV6x3d3wdXZtl3mIAnVCME//DYnMIFSe4UNTIs
WE6etjiUzmad0K3GQC99j6I3tpbLtjoDJxVb/0VOdKzMl55DDtEgerlvEuTj1ciU
YNadFvB9BxeBGk1wqMTxhtMOjsvq/h7oZ9ORHmKILwVq/o2kJ1o2MI1hgmIZj+Zh
FsIPxq20nAsTV6/lJJhjPpbcNZikSdlX8bb0XaZkaEKBrQhaewvkttxnpco8AWvn
N1GZGP2OjJf/ArDm9NCBxot5/y1wi/W+0LLQt1IPKUlpZ6rbXfA88BnDrXGYVoBM
BnwwM/Z5OXWeUxy2Ne7LMNxoBuVs44OoL9xAll4KRsOq98b9VJbvg6szNX+k5jbG
NgXRnMq3L7xxUZe4c3+dTLR0VHAFJQ6Gim+bjdIYAqN+P4hjQyf6VHGhC0kZHCfs
a6Ha2qK0GuuoO0rTJpLUZJ+sCc+DtDjuUm8PXvIpLx01nLsTcFamdi3ANsL4bUGP
4KYJLW/+BzOKEAUYoQkaefJL8Zf2zMrgLe6gsDP046wG6XL7qd1BOIMio6IjG3R/
G1PzxI/0GCGvZIPHDQcoQtb0UfT4Gx9lmEJtJHuzl9V4gFqKGh2MDV5XtTDbfjoU
0x0iVJyWvLgLE6gT6ZOn0Nl4a15J1d3SQ9G4Ws5DZR0GbGpZGqX+r5AVlKJE01Sv
+4IwxwO78d5q2qzI93xxfUCFYuBL0DH+Fc6lyC98hJuSfeYOVBwO9R/U5KjSmwHY
598dIIOq/XBeYOOUgFneFsX3P6ZtFW7mQt5+Cp7/oznRafbA6mLN5IQbbVGD1EKh
EzwJfRZClZ0rK96aarLJz1n3FgTymfcelyiGC9Afy8Yy9X1Y0qS5ixN3um/MR+1x
WYQEJS5rzN24rlilfSgPAODwomdIjTLoDk1XmAogbAQcUUu20SbfIx3xnr/j/XcH
mCKh2knKTeqru7QOOb66Sc9MkzD1+tvr0MpWNEnTJ0EaNR4bW2pAUcJ42Imu2dey
xNcOpxKsv0flw8eHT/BGXYg+Go/bqxSexxvR1dYsaGiwawKVMF7qX13ffdclhxPM
OXWFaJKujpCZUrPNKa4viPe5CrIxQNJ2C0Kzcto94ifqWq1ad03by6v/tbdc3PX2
Ruk8P3+JIjm+JX4C5Qy45ba8lgY+N+sN0v3rMg1HmFVm/T7v1QLxxleMOZCX3Nif
NGyTtIV/sZX3xHW58dasvtNqqa2LqSFMelbKQQzZuF2lrKon6heJutItj7yOdGsM
cHGf1X08WPkVMbb6d7uNbhIdFd9s1jxx/7CyrjAYoR6JQU6zhlmUWRs0LoMxtxGx
rLkEmKSj8i5cB65lzV3Bywocvo2nRN+mjWNgOWBYql7lSMikJdvY3fEkRRFq82yZ
59iP8zErMt7uBGnhlIlG6OTlogUYhVyjnFguBzrZgql662Kvt71t1Jlq7MOgKO59
Jwc1A65bQi5f0uc6/cVb0KYmGPACwNxg2D0NVMt6KjXJFRYXDSpQOQW2Bjw48G/J
YiVqjYB9Bh5Z2CvJfXxx+tB9wdDi5/pdOMXdemQkun8gnha3QtW16MRhRbs3fDOZ
+CNqOLkSHETYPS6fgiVz64BVcWhZGYxX69dusuHEJCRBkHu8WmzEhxjnZ3O9+HTo
TUDRrU2VJN57qdn9Yz8Lv7MAuH8z1C+CG+9pwhL/Gu7O9iFz+tqvuH0dpuf9D0BW
TR9tL+hGIWXmJx/lomIF0aoNenYPebfRQDA6e/WXSW+0Mfivb/qtGXL7lS41twnP
FCFLzWYURwd2HtWoqdxxcnVJbeJ77y2DeGBP5eMMftENJKLYRBnyCEclizHRL2qp
gJDKv50XMJuVAPgkcwUP2yzqlL0KMYkrWOysYP0YCXx3LN4EPZlugG7kTsQ4ZgNm
4OF4HR8pa0WJh7h+UIUPSURvSSxtWlIhuhcQ4PQL6bRk70E0uBkuw7jL8e+1rqoA
Bmr+Nu94GB6v1/DZBBKMJVvZjVFadw6JOjbM0DyuO6rfD42UX23XsHe+eD2V0+WK
aJMeCfnwrRZL6wiSvuE5U/h72GHiDDLqD6StGmFD4wuLsu7Sp6S9mUR4Tkq3YrpZ
63RvJME7nf7bQl5lbaUFY9XNl/V389Rn4CmN4+r1ciJOL3rRpCfH/E9T0hMLc8vR
EuPLLOcZPxSgN3xmVbmuSEtVcq9V3Vjhh4+WjYY+30IWcBEN+QGe8Y4/0WBlLYi4
t4gDSDuiSxH/qKL9ytX0Chy3WNrxOsYwb889kAoDLrcS/PEJG03G6CQ1nb1BSHze
/N9xV875xjhNw00gwg1d0cWA2XQ+CrzyV4BK1UlwpDTt3G5nEljhfZVZeWWFH9dN
SrqWJrcfuVFbysjnkgKp+p7ekUgaOXBD3H+a/0r6orZ0QIE6MizWb16DjJCzha2M
kWTUiZ+wLiRJbVeGmlSgLk89k/Dn4/5yxxWBbQdC+HA6HT6noK/GyJ3sB2WO11y3
yAg19oFfOIOoQVM7wFHsPMWW2p8BdiOkP4aFhlnx6zITU5cVnDVzHNXOc9s4EyOC
Ax7E0k6dkOcGJ1mWTgMu0Ms953n78srvt7wS+dLdNGiOuXQ1+xh0RQmGMLYzfyrs
jncptlKVb4EzlfoRl//otkwXA5HxAgl0Zojc3n/kQDK+DBhpPsq152+dEVOvhX5r
GThbjms1fqcXNSBtlpMSJRpC/EspTxxIi+DPxwArKMycHLxAwO8fkqxdIJS9VcxU
8FNhtIAJIOuZ5Q0Ck7TDhQQl5e1oliZsNoJMISnkU7speo67XjSsGeX0rBEN71t2
0L6tjg8ATn5wdVb4sQ9CYOt7YW5WOxsYZh0S5wHqSgAOcYoliUed6odUf+3uHgly
BypzvJD1k5mh2D/dQwB0+gE0tltLqkaZbA6rRXgIF4aJpTznthfAlxEF9Dq4qB17
2iPTA4Q0AVHEZuF61pIRb+VmxL9ETn9JvZEmyvF08yIIAs+XHm+Kd0MZgaV4mArq
iGGP6LAArIT6m1BwC0rbFClWVFVz1aDxZqOQUS7xlOeHhrVZYSCFalpMmu8YrW/n
xtFh5GxgMN91ncysP6i4R6RBJkfaXYue0KQ3lFzl+XS3yB5YDsy8PYPpPaO0OZJl
blU+R46pd3v2t3i4Q49BPVV0FBO25CwqTbmFHk+BrgGi9B+0BiKFJv1i77xk39jG
yTWHteYHzIGxTbkH0z0Waw09l8uZJtBUif+iE8dwtPZmCt08zoMfutxoWQE5aDP7
30xis4CkmnftEPWXRMU/ZIb3jKqSLwkpVv35Y0pKvY+Ck/dWN2gQNWH3IqXzucXZ
GiFUleyrCL+yK4sEMwXJBlJw8TCA2LBW03bpGWgPZnQW7D9sjp1HyaYuViycw4g3
drN/0MvWLzoxmoTk0oxGgIW9Oy3BQjKLQl/qgT5ZZN87O9wyGRgO4mipOxJMkiaF
nneb0r5ccBtKF6ez66+6IRA2ZymUEy7KX3vm/D/QXiSn+c513r1IKnBuhRz5bmUY
17aJGS8aeccnrbiu5YHACTETngZLfZyTKenrU10CXz8CHyYbbCbSgv7PHHaX1jrm
EOkO8a/LtPA7UvDenIZp+3Bxkvwommxob7bxdW6wQ+P3ZZ6WlEPfuHMwCjARvSZU
2kSYnAQwYTDLLLuuWBondoa6+VUjABNK4APuUmSbf47VSiwQB8uX930aiduY57N2
rJ4saag5xTTxLBYAkWIK5QlVytPx0txRwCSJ7R4E8v76qAV5gMcwCR+ZS8+XBLXG
sw6UtXJYpF9nAakCQxyKA90sCtUP9Vq2IjVOCvgzI/+gL7MX4Ly3X8tskyQ5nL3Q
mZGTsxkR8Kw8sxnKVnIRm3CapSh+iX54yH313BI2Yl93vqc2E6Hz5DW6wPO7ovD9
m5blGJFZxG1tdt4PWOhMpXSOZXL3aF7PgeRLc9Oxk1KTvF33DtKsu3QmdAtKP51V
ck6at8OVCt8cIrzeeUF1q4Xp6JxxhhdDalw8miI3sFni+NiFNuXBasn8LV7grxxs
nr1oHopWc5OKtW7xGS7dibuMr4Eb7Ow8HeT5/gbvCFZjESJALVVOBPbdIneQ+dJ0
fr3hQLkXIfcg6ZdMv0I0vq/sxkb440R7cNjgwfUWRul2ZzaWlF5SDogc39GOH8sK
MNQMyMrqbrhODkNwXWecp2GcMC3tEfZLR8Z3h9jpXgMqHJChDQuag0lz7sBC9ugB
lMrP1VBVEcFDblgdbkR1y9h9ce02wL8MLOIkxhNnIlM/ZSwfL9cP7XswrldHe3TJ
X6i87ul25e1atxw15gunM3nWQhDVF4358kQjKolZVE5wtt9Z6o6v016DfSxuIWZp
hYFpmFEIO3S69at5GofU96eTPQfvwp4Se3DWabJo8U1U97FTVU5t8xHg9o6lA32t
t/2N/YHDzFymrZ3asY4/QxdeC/IBzs4OFHdEDUixVbvA9WiziCF0Dv2hPmFMQHs9
R0F/RxUx7stIJsqTUmlQFCqysacHp8kI/4aryDf7UJg5/umEHNMns3PKNWqwN1JB
Z4EnCAAKF9UizueIcExUac4OH6miL+M02hrqiGDI7U8n4ep02+JsJTQKhSsRJyx4
LcgcLGiTJPayFwo5mmaLf5hZC+Z9YubOIW4GAw/73AWnC9jhqH5zYl0YhvwrRWPQ
cYfAWSQ8amyxyiipOBl2zNncPk57gHZYdC3IqWpBusicv0EpaFK9IMgWilBLnm11
YmpmXPlIERNjWWWjCMB8HELNVqccmS1MdRpePv9tSdYRj1j0+q2+EpR5jGPq080u
wNB6L4wncOonTASyaHCB5c5OiR3ik5ZbcCe/7+dM3MUWOLscax0/tZMKUJEoQZbs
C9LLRoTuToXnwmoPs/CE+/mOaS2XSu/6heEX7/xLNW3LfhnOW5WsMzE4MzJLF8/p
KZwuBBvTca3Ue/x5+axEhxg5qXsryohSYJP7qak4bzMPepkEA71Kn0OejZFMdTmp
Fhqf2+dpCat3uG77+iQYZd8iC8mgC8T6HZFOhhNFOePHkbsKcVYtd79QKchL/8A0
5mOsJsJ8u4OxZFBbRYEZtdZKMUXDtRA7oLoLhViYsc+x5FNLZqIBZmOFy6dEcg/g
i3QptvtxGupvEVEdJbY2KTz3uFCd5Z7obQ96G5iJ582JW9M1nxUiyWXGwShWC1VG
tPLD5SHJsC3jy4OQekm3aqQkjwAwB68V5/aKiX4FK+iqdGI167UABi0GpcVS3fTJ
fJ41r1EMM+QqpXXWAfYNhljMPVUmLQxZSdrNLUW9CsNcvgyYaDTO2Bf6nqlkOTU/
sKtWY3opW1cEctxhPDB6olzDNHTb2vECmcigtIH299seh0vS5ER+rDTjtkuE1dNP
xuSMFv1RWltlRtI2rjSsoSjXLjR7lNCci8mp7+tuv1pJmJqu0IWzfsTPSofN076k
hiELpuwc9jkZwvcG1wnnPxjXfhWYvGMMEiz60Cbtwj2VEJaJv/UUXi9Cfy1dsPeF
LFJf159SVXpZd6HeHV/JNKFKpr6AHLCTSqVQI1CkpG6q9gf7eCrR65OWL+5ncri1
j0jscqFTDbbjyqu1pBkyXGOgiTCkY6G40nKAgtZm7ob0suddlWJN74TRTKF9p/HT
ACbDrYPeU1bLsaMrx4grf50NL5xo555r3QCnsaEz2eUfTmvzHVJr4EvxxpTGS3V0
f3p1zw4BLVmVTMB70SnhmSsucVobIerAROscddl/NL7UDMn1Eg3Mq4/to9ZILj6k
Tb8qLP2/ovMwEmKD8nwqvNLM2lIfhNI5qNzt5duTypSH1pBmxidvizeRnVdpUkDn
9Ro9IzzDepGTTs/5VFeBs+pok62N0myZW9ejqwfksNbIee9GUiWtXUDmz3EFwFAp
8c1fkR9x+yS33+geBaN1Ul3r0vIcWWvA5m0jtWLBG01xBRSV3WvL7+iAbBJaMBCN
j1nhsZsL91gZ6H51Tv55dbrdYvBFd3/AuhD+y7V3Cmd/t2cw5pJ1/xwE2CHjEfIU
xkl0Zkh4B1YyABGyxKBXPcjvViPyIPnsSaWKok6O/UFFXFGGcdgeqIAHoqC5EM1n
k6zvubT0NcrHW+oHcPOyIy4pDzHoqMTAfoIAcMHuMrloQOr7ZHGrJRaYdyWLDsry
Aftk1L/51OkuwsjLxqwc9Vxkli2ruKgtKOnRDjzu0hQMv63fkZqqRsB7NWPMzVYe
NljsLapgUwz+B+veHDWWbify7wBoxvohvTZkW5wsHcHbqC3pEr1WMN2hZ1bInZLm
0VwIDS0ZmOp0vE8gM0kBnFXGPsHEdbt8+lTBpA7yZO1wHTbm42QemY/rDz3udm/7
IFtv9bqgELc7/O6Nb2O5cMA8ED5tAXQR5p9T9SEwq1D5SVuBrO/wYAOXiO8VR+wI
iNBri4ckPccihfz3DIscpTMuh3su7qWDttmzIZtg850d2E9Cy9sHq4XK/Q9auiqf
ZlVZKJlGi+b9cUUXuEDwl2a9PDoQb/16cruWMUVnEiceADwD6ORy+faSDyVU7LnO
N/83HQWOXpmg5lew5EhFv2u3HTVxxt2bqGzlMcDhlHSWgvxW4zeTFsbhIN5ApiXt
aDnjOcUsIrX+yloImSIs/5HARzss49vzfUq9tqUCGS+4pIihLR3cXK/TMVBHDseo
CVgCer7bNgBlHxXPHF9fchR+zYnKlDmmJlOp0PsgRGObZavnTBFKX0QQ23NU/SfI
Psd9TX52h0vtfq589QGsgYRoCxiT5+7UE7AlYLHePM5x+1QTbEtSN0MRW3t/rWUl
prMazP1sxIgRxA6FRQCB+omgmxudqTXSIe0piEfLYMcexyIW4ZObt7hrZJtd/BP/
HIoh1CluJTvFa/8bsL2ZKA1R1oZUnXVk4weDnzcEy+uNVmCw7DQVO3lmnheOv+be
STh3wHibBxrZ971YGTfvhjJkeC/LFjun85YYS9ctm5VTpD91sccvQKQJC/imJCIo
zjogKZOAOn1pImvxk/OUvjbt18d/vI9W0VjvZwtF8qXs86K/mhq0P7AYI4GRybe/
4Bj54zMnRwK9E64lbPV3B7pD91E8sK83HjaOIawdmrlTMW66azLN/y4Hiu7g+ih4
CKL6iRtS86+d68Y0bwisXUrDpJlAJ0jBgiTZAriUN03NGLfxOrdBED9meMXuOnd0
aVUR+Z1kEANBchn7b5RQXmp+rT00tF+U/uC7ILucBXBpn7wVDdz5UtRepzDYLOoQ
tA16IIDFVH9Hx4m4X+JeaOIL1qKzPDigN49XX9kBlkRnIPwa2btO2WKu4J/ye0OC
yWLF7El9T4CQUa7cspglV1S6Ue+j6yG3sgQ+OSF0xQBYQTaXuU2SUi6hESugfaB6
Lko34JRmlRejjK/A4bWNta9ladxKFc9GbSxiPgOlBVU/pfhV4RdsHJR/sT10+3o5
kVjSsbBDce8lUxD1pmpg/T+BQNlkAKTAjrI3/n0vWOKADeE6QaJlX6YiY1Bx/bm/
hE/M4qMydm5NLv16S+AVm3aF9mpBzEpsVau5s6IAoO3J7pe2kWx/W3h1cCLBxFMd
GoeDWmrJCPf9uDZaFeZrKdmrisSnfJ1qreZ5Cyi4a8uLEEpWcjei0lT6RRgF/0lQ
u7fKghTkJYehipSlYjtqxWhrBi82a0/Ds5f7hMe8dhDqkI0i4lZkVQm5auN9J+JZ
BY8/9CqoHLFMmQ+3/vumK0NJi8ZMi9A1x9qLl7IvFNiy+IEl65pZbBnelinNVRxJ
XgQQKZLh1GmDKPswBpk+AXupmhKZ5GIMsV4ZthWQWb0XZIcTX162sYD36/AmIwX6
vP8xuCiYsEI+ITqjB8we0oVLiViwvBfFo25AVYspxsEXtWcumuuGoa25Gs5jn+8q
QBqgiI5s1GnFoscH4WCmAicGnTbh2Hipg+Ni/wfDW+HXz30tGnMAHaPhqdjxGt+H
SO7WnrE1wDcNkO4Clry6lgDlJo7jIBcLUnyhSBFfUbeHUljAE9VQsMv2C7Mg1tl9
BrTuvF+LllQBss1iICTjvWuiGEniX/ku3jrgtB9ex7kMxhd62EzTvgWuP8YvRTB2
d8LzhXHvO4UUCIZ3pXdcp1N6RS4jy+DqeYXv+SN1SIXEvuGgcgGIwQOuWt6uck2t
EIim1L6rDtTZ8eo8OxlmpBiIsg/FJ6EftvW8mna75PTCKpwPgHSYRp0DztXbJlu4
nw2+szvYaldypnEFJON9EuWyWXbsyyIsfCLmrnCYAaVpt087kAllgYzvpB8DTySJ
kmvazapow7HS3UbT/L1lhD7pcnw+vYpzFXZFsnPPHoPVwygyKQIe3n5gSfKt5W6g
k6kA3qKtY+3S/xenxU9GCwVSRk00vvCYZ+kJZ6xA+psEEMcC/t0fXD2MrYp7ORpO
Vltc0gUwmGgR9mcCEIquLEHQ9BM7mm/THtnzIGQ314YQ3s/kDc5Y9W4ppfmFn0bm
bI7K47sMI1BVy/OS0iwisFcp3541idoFglX1JeskOJir1EbFcuAfTg8PZr8tHtl4
pfEElOcIVUvgHEgFZBZnB5NGsWML6nTM0JBMB+Brx0+bHeHjhwnZVaWn/irZnXcj
D8tTjigoUzxNUz1JEms4hZOgAE4RQBQ9gJ2wbueh8iVE18OOjlyE3a3Fo6mtRR65
H9ZLL2moaUdt0Jd6sjZhx2vBTW84sFH0XE8NBR4tcd6p/vW/6jjNsERC2u11XRE5
5WLkSAYOIDXv7ieg7MNZaz04rxbJvJwXtGx0ZT9AjV74AV8JgPO2sCqKATiBAeaW
61atmnq84kXQrde/3K+/qO8RGmt6xPIJFUxfZ+ziHf86mbJfILiAzWFJXNW7/tBj
rWXoibkrqukOLS1LLOeCGRTmnVCMjSNU8GxuiAgKfNq0H4/i8kqilVJpf5RxTjPo
6n8MSwbtSHMdV4V7n106hJ7ggVmGClXqNvB0FlG7n1toaoN8Jlg50UJcAgewmSay
dKx67RKw5cvOEYjciij+m1uEuRfe1PYlffm1PrIZTGnaRXFLTu1fTx8OqFtPotPD
NmmaLcD86N0KeAJfC9ufs7QGVZREAl4ZlhpEe+wtfS8EUQ9EUKPDaZeG/vWlE4O9
dPh/j6s/4s/aPvOHgKuRImo4SeZv4uNuK2jI9fDZH0/H6V1L1Edf0ivg1wv5KWCt
26kgcjnKOviq4446gdm8H3sAMu4V9M0paSSemviuVh3VFSn9FpeUsJcDpEVtgkdu
YVhlTbfiPdOzLpxx6R/7nutrhrx84QeSa6VDPEpF7rqzJxlPxdpO3O3O5J5qVJHb
8B1O8ybL5ByungtTTfqyRBm5/GRnIPGM+zr9lZboxjCc1MPC/8UzBH52S2G9Qo07
PN0TZ3V15LBanqEokKUJPUHgWAV7UKkuD2r17F5078PpBki/aDcjTr9BCH1jxpk2
pQJBWmNoco4XjtVqLJfGNtyF9NkDTDU7Rn5o3CHv4SHTtc3fWQzU/lJ7lk0WnC5V
HnJaYY6irNG2xHBDDl/Amh0XQAlV/icsNZk1rIUF9eBZShV1hYNdJzmzNC2yWhjL
u9tH6UcCnCGcfb+ahfBbb0slIKQ2Armpj5BJw3zT9wX6TtokndzCVi1ioPFEb1i4
b5yNr+6V7tMdcFr/BcTb5/LBuFTFaXo1rEU1SdzLmav4/NrZPxVO7Al4BI+IETFl
rrplStwFQrSMwBRPR67vZ9zWGrSjPJVFKIDHbwvEvGaK1BJxWlWBkI+C6vCdi1gm
5/wKy3OJhZlhbmSetsCTzSCyy9KbFZVQ8oTyhoJULfD39ia3mmyNajlDen1qB7oT
I0HimmUFxns8bvpQpPiXOyjodgikTcqU+d6YpoSdPPEhHE1A5Z9kjbdGR1KJOwyT
QQsQAZl7UDed6GMRavA/oXI3cBX635s6X/YB1vsC43WOvWvQSXmCdMZV1YGXMOLI
GE3J0VwcA72W8JkvJJB/tDdA32Sv4+8L14xWZyAXCErIIbNEv/ViNF4rj0X/zUMP
X/QgZwHvKtYJVvQaztcPXKO9sV2KF5Qi0MbTVXIpKTWHL5apFdIBKIvWl5jE+hJU
+8AavhVmTfrm9Fy9I0UEQQeSnjHJHBIGJ6lsnJYN4x/PhrGfSkkT/9Gj+i9tRA+W
PoFyjPNKq8sWPbkPhEBmrPBxRYh5jEGR8Wxm6b7S0urvW0YR1qps65dGmhX8nl/m
uu69lx+5qShh17bgiaNGtmvN4Ut+UOBr+rDI/U4B/zWj5kDEX4fPW4YQ+hT14/Ar
sujgVvIHMvV39rExBBwpN0a+DR+NqCTzT/F+o4JsbWl6JeQ3Z8tQx6xQ7zAHfBwb
ZttggtVzL2oOE7zWrhLcLwA6AZqKEr6gALTQBVdOFsw+PuSMPfWSQnz3cQkygmOJ
JI01QfbL64+63E63/Azx0dESzIpFP5lmn4D318qW5TQ3Ct9iZ6ldC7fIBzHdGmEo
nVDbGsZxNqSoYJ5sTc6xi0fKsQQTN1JKDodZIm1NAZBYj+uaSz3zi5JGUI93/s7f
9hjsbOJSNo11nztaW2IRyZPPELx7+MaUyyw1uiv1SvfJKDFvDlpHJuJjG1iy2xgM
TFBwSmsQopVP6WwwH6E95s1CnzUsDE0SU5V78lUBrQ7tVsDN14udifuGo+ATJnKz
TzOu6ZANafslEGEF5BAI+DbY9VOCbe7xSEuvZW208npmLa7EfbBA6unY+Ph7n5eE
CdbZbsVgCBarxIi7IjnsNOkGRL4MhPpOj6eP9Rgrt+vWujKwznwb6UptQC+4jJfg
EZ7H/a6RTXqqFgFIkmKRMBOAcNZPPf94V6AAIzSiz3Q/2jdpkv/dlg/AiUFVpOXe
bu06JrW1l9di4KqEFKeA0YT3SiVTf94dlIwLLDLS3EnUHn41TjRD9jQw0XyGkilV
Rs9OOcDocZSzlRoPiZ0S/L2gP0DZJX5T6sUyKZJnW+XiPFTY0ziQBZOG47wvDhJi
PNtFKTQk7WfRaIH7BPp3wfN4gGB/rZijvXSjizv7FY0g9WdnbjKd6607eXUCLJyH
GAfY0mYSpMJMGtLgqDv1OEOuHe0VJanabvqIuYUMFzkf02u5h1dRtsGfK70kJHHh
P3m0/qhUBY71at/yFqVbte8/Md/DpN21WtvrrBhpwt9LgSgsJvtxPfVAyhb56eXd
cmHSzcmNvTEcmvnwUxXXaohdSb4L8PD1OGZcK1JPw2ZsBrBXt1y1G2ZEAvuHxBh6
fzkhbi0CDx7x0aNwGkVLUaybR3y8d9aqVARvxDrcKp/nSY+bDdjhU3DaerUoIuNz
Bx1IZqnKoj7lVZO1ht77UmIpV/LCKla69G/f08ZCAnuq5Khrpfk9Do4Y1As1srsa
8RzibZkSdEF7eI9sC+DnX3NOGTwnUgXwl5CVIbD0q+Hq3mzc27DR2Mq5aeJ1btwz
L+AZRnX722L5rnBwlaYUFN2Nmvx+crwCuixioaq4qRYjVMIXpdscjeovJe3lgs/b
v94PxTklDHAHZbqPKpk1SY+GKSTZrayeOg6Cl87xS9TO4wIkwaNjJFtRoJN6xQoY
sATd5cZJAI/UanRg3Zc86SyGOeOs25DFM+KIOinVy+Zm7FGD7ro/wnJPP8VHBiC6
pGNq6xnDzfyIdodFlRj+m0cq9J9v1DqA+nfBU1vtj8hF/v7EaybFlpjPJlTzKxch
+sBirwUCEIsQUBvOr2iTuqrkbMM9F7FjX5yZjOZUTM2FV+QsJlD+4H2ooyRhNqaG
t5iYw/o/CYg/muL9cfbgTim3ObeCsYgHqTQK9TuyWX0gRs0kvW6SHPqohooY2p0d
sKJsJDEn3ndyRSOWNk4f8lNl5q1yWsba0oBjbRQk3ChTQGvU8HHGqDGmUUvlQNGo
Dg/dLw7si9dp08SMpdeLSf0C4eOew6Qt6CKms0g/4/8bNf8EqqmSaAyxyaPAus81
P9fnuZ0EVMQIN9MSbTQVED/zej1i3oEbKNJtoQ4jl2GBRZQhz4Tb4w5QlEj47VKZ
TJ5nsHkzkqXA50JoUhgrPu9zj22G7NRR4WKXtEesnZ6YAPUm2l+ghWOO7Hlwq5Re
2cfSPGnNlrgki7fdIxngKRxbL23ps1ZFAZMkMIWFUyeZe/Jx8YErN7woXik3kK77
3J53j6f9MWKUCmVt3C2fFKrrotgHZRqm8VJqmLm5ObTYtkwUn1TODQYjp2LcRosO
HvXP3Qy61UwVg+FiHLpecz5m3uAV/OUIYsscpIGqyZwXsYdX+1ldwX1vEbzjwCos
bL15gyI3gmkiOvXhwCDxMbzAcYeUYEIU6IWIXbXA2P2HkFlLvuPnw3qyLlvr7GwR
w6GKz3ljEDBYi9z9a9ZB7zfOIjnDEjhzIPnVV7q5IC1w6yEF77Eez6WIxB1DOrD6
V2YpU0gpUnAbJtOoqUbKArfJhvEoDfTskn84bh3rwKBzJS0GQCj4Bn3/+oXN+vJ5
ERZ3sYgqnqx7ZMGyzWr95QObcJ+unLsy2/Kz6rrRw5zojJ+/KkSRpT9anSs0g2yp
WsyWQ6PYfyc6L+oWgi2F+wQDmd0771GO+TLgLH4ArMv7tYelHwKoNvodJk4VNIu3
VAunOrA+z1uAZQWywUkzt7aX0i9tb/T3q6nsVjIWYXR7LhxGza93aWzuNd7aDNQk
lJxELwKC0lYcv10n61ohh9Z5WLN95pHefKQCAL34Z9AShbetIF7rKBHWo/PC7+sy
BtflI/twgJWadxryPz2CdPzcIQtThvT0zaGgxVl51RwvHmZzhJUxNqNVRiO0g0Z2
BbrbKjuH2gpx4hkRP6jXyhiWP/Txptr3XO5vy8cYtYoq2WryNKj0qq0LO2Nb5u2z
TAvmGODqEsfOE/t1+4Px2f+6CDbbqfc12p8nSkxRxjl88Uf2BrAXONatfmLsYscL
YloX8FDpSU3Rpem4UsuY9bM5n198XWc881SAs6yr2Ida2iN6p6NhNvkD1VCx2xRH
UVyx/5GXUU5NEihyOTugLh2dw5YZWUAaeR2UTnqL792H7ol+rAXQRY6iLZ65iOAL
/kzAiAdlIzARfGeTewr9SxV6E5l0rbmkRkxL+q7nJz0b0IWgLX5TjbC0v6bUCl3E
8C8CFRXe6qLZrpMmL5XfcreWem6yOFlqBp5qaAlBr//UrAPvVCub+xk1raCprCFi
CtpFeW1AOLVzg8ZXMy1gBc5XrOlwcuVZ/TtHA/TdOTmy1HS9VxP1KjaMa6tK7tIk
9cCP8d3M4T1A2xETgkzDObhq1UpSLcMnIQZVrGDHup8HR0kVOKXVfDCKeAg2REHh
EVlMqJ5uXf6NUXXzR7lYVEfcc0+QfGDN4AtMGqUJERoZ6rfzgMk3spNQb5LnP9vt
JzHiNIsBbWgS6Plj0TpYh28nLHjvoxIy+0qGM4OW9F8tYC4P/5EIOm7XGQ/CFeE8
4KrSNdb3l/QUtRVXdhujxtmf9dtFwxrfnjh6zGfj6hiZjzKndfdaaSmBi9Dq0t2q
2RJJ8h+/ZfPq2sU7y9/GqIGSnMTjCLfK0LuwDTTcaffIMVqRP2EMFT99q5BKpFpG
kmA9QM8TjwEyhUKNbo0UGrFQtuH3CWrG+4vigi6nlVBdhKSl3zg9qTJba9rtM8OX
6zgYesyyWxDl+lqaJVoud/PxpA7fSHhN2qvvii248TH+raJyo6YXgqCU0lWPUIS+
ZhUPeoMuy4qXMSS57IQo5GZzNVDa7pDFMtTcNLPWRCN9RIoSuvFH8F8c38k+M791
3536PsfR8d7KECVcANxfp0KCnIYOtyLpXq1F5gCjVlolb20dkPCnyQphSNMa2bgs
Fq8F3172d2hEDta8jV7mR/s47aMtXilQj4aIAhgOUkpR0gyK2Pse8I+nCmardN/q
oagcDJCP1bUW9zQkbyr9EmroXByL1R+AvPdSox0FKbsv59WynbKHshPy8zR5X+7N
r9UJIYwA6cD8RnjbFDQ/TlcZbdDC/q6NYOGSEPTmgeVIDdoEXjVdQuoXMAs5ciZ1
EzR1NIqefh34ilLFp5udQB3V3GexN6hfixkAQDly0CJaZUxslcDEpzHdQ+uxNeio
WsEdt1InMOIbnCA88Rwq7119/3WltF5RtwvdZFC59wGx9d20Drdwpsm9XTQ99qOO
B8uOVVt8aqwRdvU9SFSjoc0Nfr2TfAiOxZ88O/mSTUKlMqZDA6MfVUpXwi83KkxN
jfmqs4OBTs10W55ZxuRLkkoiS+ay0NfFJS03pyaXohZx420OMzkDxLlkYJi3j4d/
wmPfp1gZhd0peRQDfUocdsIGoGvTxgQ6uOWPuaigVa/pf9am7rKqLZVW+FqKJcmd
Nf8KvIXCv5gtY2Gai6pJCwKOd520PCfTJ537z/xuQ8n2UJdw2LtXfskoBb3rn6uW
mHo4gwzIf5sjbHytnnpN2EVxuOExJaGrhvpB0us+bZXswn/PL4kDthohv6kCU1gx
sUEPLUbdrnx5NcvAnswxGIfUaMuAixN8Y/bPBdFR9nmP42mRoJBeoF32G3TVmQUQ
RZH7LZMUj5mtuVWtnvk20jQfTzbELpaNVC1JEzDfic+JtupCG7gAOP5rOJdVkghg
BpSCcflrzEYptgmbKEkpqaRY2urMaIbMTEkTVl4qs1iHvihFuFvtrI/jwHHVJHmi
n2WeZzqiZLzBGgTBthfMJgJz0X0erbrYcdeBW8pQm8l2aTWMC1ALNtwOyml2CDd6
pHXQmG4oYZ7YOh8vLRimcHwUhbKTNZY1/SVRlyQTwkHc5Nz3D3w0fdjv7WYUJpjd
3gRf+5sWnJkSQ9+YQy3BlD1Efq8AmE35E5lO0nHOMNYP/8eZ9KBWzUAKb2JMW7WO
WBjbTCXYHmjD7GT+rPETg1kgZ39ze96jOTUwt30LRIRH+4WS1ggUoiDzT437Buk1
r4FzH8T2edqsA3CKL0EYW+KwpfzZx1RvJ7v0CXqjKZzYDawONCy9OzBjYqtkjmNz
oXzPiXc9twx7xDX520QwHEfYYok30Tnk1y1boJUg4S2/vck1X2E6BSEL0pY/LVbh
uTNU1NurDmqp/ZZG6oCDkosVdM2RBsIoM8rq/kZ1Hzw5GlBcC5WuDmXZYV8f+8gr
z6tIYljs+81+i+4I/rWEFyvbMvxGXo9JQJYzLqC1CIkOsJQXBTb0WVvKO2FPZ1qo
hjvOlFitzbLEN6amsBbFvsIDsVNlYTBXSOAemh8l5mxkC5xdZ1fsC46V3fplVgJK
iJozfa1quIpaBuPuLp/C8tUD2oXBrQsg4yKsLkiPP7Glf5hGpL/9xoM21UGHWktm
3+5gwoW9SP/A0pLe1Pk1yFQOZvqErgkS9vznyiWp6TWqFuW4qDaN310ApdVs8dnH
xyBJkfTodlTpzDZO54dDnq/g1NlylI5ECY97tnIm6FJTW4Xm24QHx0yykEq+MTxy
oc973/MQQUy9gAopBZuMZpqKPoSyeITN0hwTRYGRjY2Z3RBnnCmMguThs6Z8sSUD
8W+dQP99/KSDR32muocyKQTIzUDyj8O/jVvNshMyQdKC7niOz27vpiP1WOO03nVd
RtHiPBAvNO6RUHRTeO1RkosigE/0xPFIYT87UrxxPo27XszwQ06qkiFtudnb17cF
olAlan9T+EUE+djU++4ChH92u6TNolIICFeyYKf4V+m00EspiTWEYaFwWV9tRIc0
c9T3TzVIGKC0/gjRbxPaNExh7Srp0erVbx4LZQEgLUCodIEdN55SWZwEQjwtJv41
09qQ1cTzlDA/f1J0FLBVz9L1vLk2/aGGfO1Jl+h+jlb+1tz5YKRVz4fdKXJW9zYt
EPbBt03ulaw7Qfp6lmuvQQRhvSXiJ2tBzGg2cjscbqsMlb+lbqYL6yK9jQK3zy/k
cWwjUzGTK1PfZt+hl/9sbxPXZIGuUpkNwxHYrRZGhGCqv2JM8dGB6+CrQ107+Hid
oNXPBVPm5ls2w7DAjtMZMWu7WD+pP4sGTz7WFONBRWYWkGxDGW2M4FIzJ8p44Di4
+iFZ6NJQsHui2jzQ8YtXk5ooJKpOa8OmjfgeI+5yBklb+OzZatxV48XHepYTEvFR
SykQ/lpqJFbH7jQEEzI1+sSI6FLSBWwDVTKZUbuCsFF/ALYb4EFXnouAw23aIeyS
dQ1q+DKqdZByjv2hBVoW/MiY9jwiax03U35UuQqfmI0w/AvXXKQVCKCfHiW+PVxQ
f3zMW6xCEqojkj4/YTdo0iRDf8P9XS67b/AbDiPpzIRjb1XNwmEZTF8ZWfKvh8Yf
eiO9ehFQhUmr6jify6MqwVdoPiyt0PpfbL7Cs8Q98igsw/RFlx1RIaYXD8yypPZt
PbaRuEFYm+IUtkpbkDFVjBCIUcdtGWNXd/0OfzMxnZYcy8txXXsL/KN8Pr292x0b
ggtsMZ447lkg5+7Qy53wL1RdM+s9TUTZk5uHvU05MLO2oPtVH7sOrBl66evjHOu2
VIDAFFiGO5CnfYdNGTxRs2dBu6Q/rMHy1Gx1EHCJDLvvkc59JD48MgzKrAqigVFH
GnAJcraQXOoOpLlLrXBK8sHMJNn1RChtrkEpG+/8mUb69SsOYK0vNPN9PadHQTwb
j2awdZYScS3ip8EZp69FdavPJFBp+SJyyCnOl8sSE2mH6MYEsiYzz7mVndiKoY2L
a6uOxkTNfc2npRlxFAkngsBAwz/o2AHsZ21c0u8LLh2XmUNRefQjCE3xPvsKpFEq
JYrmDpa7nRpKkI8v0sDuZwufZu7y9In5Rc7jnvu2QsCdZurTuXfrtPaTpEikRGQW
NoQj9DOP5LnXxuiZtyCZaqabvxXHdFUX1uB8xc8iqNen+kIat7oz9PPhVOKzw29N
451EwKcA9AsoeEg2voNgqWUlLb3as+QU7aRqv9qA72KnN1igxWHt3nxRrTexqLw7
9C1mH3af2p+JE4IU/ffl1UComeebiKdaKb7LtmxU4QHExfDkjyk45w2xxQneu0VU
CGI5fO+RjLxDb8Pj/u/H2VGVR7cGwA/Sdu8K7UvbcA1ozyLlZWXISAOmMQdxAVUK
7cfEm9a6IVSUNgot6bjKKYbLTei6mj2PmM6gNjUrIZDRhK3JUDaIWZNREEn/blik
zBCot1/ts8Da4W+DWTqV/but2vXvjzjArSVTZcR2ExOzEW6epR1C4cdwOZZv1nGA
+bKQHqVJWAjJ8aXU4ovGupWIGHDJHuTpmQd1pzGeOtr+g3XBh+1F6EmBpJcaM3ax
fF9gmdaqHp61UthSK6lpXt89MI7105Y4I11NjWZfM4PV5wkpfNa5wl9sdIpDD5Fl
hZh4UhRze9O7LfamTG01ctfJ9cI+JErh/7dV8e7+aFyIijJWc1qepn0iM7i8/ZEu
/fAn6e0eOUEUkOw3NmN2x0XT2kWsF/CxYC2uOkBD0rnXYJqmVwkIUsc8+WrjsPoD
dvCX6ZqNZ58SzEGEJBao0RLymGHLka9VxOi2lXVLs9frrD71UfBIYHvluL67wKTy
/ZdIGki2l2Bl8GHcimpfzsn3y58HksXzaOphUtElRqvEacRZgvf0pLCno39Xrn0j
YEgYS6Tip7iAUP1ifafesywtV8tJ0JkBkLJHvP0vCEJOUOJSyzyWP8A4Gr0/wir9
DvWQq+CFobAhxtC2qNDVhxH6uLHKs7fe6hDqodmbYI4xh3ifJ8/zoj3s3RlzxVzv
rhI/2yrbJgRyE4xHtwMfXWQag53UgejS/jHgkDnipzepbTNn9rbXRaLmXYmv7vFe
AM465iAvxPDiCgHyH3v5050UeB9g60ZxhJ6TsB7DKHQrO92KWC2ZqbtkS4qDZ6Yy
q/uC6rhg/c+/8wMzuCHRhR8ceu66Hzk2Y9lJrCjoiiOeJt6lsnGCRvCv7Jc0NZ6o
F7tsMBzKUcsGgKyFay8QJYjF8hRFNl8Z0rehStz3MvimvhvOKmVACqBxN8f9JOfK
8FtYGn7e2lK0DEnJa3UreWzqyBXsYZh4dEbbBAzYSTBzdIZfCiiMr3JTTAmObBMK
KIKiENz30UZ06GF3Zc42sDXHmZN/d/2aBnQxkwoMetiR8dvPHvaRk5Fc+TYMtvVH
U3UHh+iRsBLbtvJWexJwaRZXtU26btGJWPSstwUUM8jGHRDGS8glGNV04rKwtNHl
ANM7QfcbQ8RlgibYKa7zVAfb3mabcPkwb2K+M3H7/OHckj8xCXE7uZCsnQnxAJaU
IG1dYwh36wSoXkJ8ZEoAaFW3Qe6c+fNebRxik5gQLyH6Dr9QMpb2Q2uN+mzZVXxm
oo2Jy8IZAFkmuqvS13CI7iw4i8dZ6ejpJhzGNFnZo9OAvay9o9/7w9gwGqjaVQLj
9+Gx9tzsqDeh2hHC2uSNzkaz7Dblf3E3AG9jd/EE+PjXZ9w5D9mlVVL1L1Cn+aLY
6GpPumbLq5ijCem4v/d6Vp/qYNB3sW31Wt+4wTFeA3Mc3+9KL5T17zTBPtq8k3b4
zmUjpu1ZWxAcR/qKwhSbFVFKTHt+rkChvLOP5Q+JnjljvlLPf1kVEt62C5feTTkI
fQvW5Dt6EQzvSmHumkensxO8gxkPnKCWKBR9FcZKyxduC4Gws2Be/cOAnlJ13DTn
jKoQeDNOnw3jbQ0JFlM1oY9tztzjsXZqadK8K45RChMit6PS96L+KUy3I0ngoKRj
OCJNg6zrQxXXEbE0L9PRYU9IvobL7LPOuuEPCVi6GjKlETujEuRTPs9lPnR0V4bT
qxVtx7jVHsYNe39/v+ziKzv4tpBYk+iFWNYJEkK7xZhk0XmH6aDzcStaMn7rbnNU
c6kqHd0Dupdzi2o2crdBaQn9SyTCcbt+B6DuOsEtwa8bZHdzspxYjj4KXE2F37Wj
agZ6qNZtoWtI87WId9DXDi8Ejdop77m4KT0Idnl8k7pbErJQOXHCHtFxtSpqCWNs
lkeVb4cPdWR8zBhXx/gTUsi1f62fbU9k2MIyE8f98l/JHrkWoCumSgVRZ+KW9enE
XI15EJ1f1UJbgumdWJnOeRyRg5jBVpucC6FVWboCTN9AiuSBG6ZdP6LPZjqQvYKO
c27xyEDI2bwLAt4TM1FW4pimql9G/zVYSRLoEbsgEi6M69Hwt3MWDS24n5t+FSZw
9YOnb/SUzlUPWvtey6qikbbFJ6MGBf6ZNn/ttnRnmiG7R5QJA7iASkuYPammQRaj
ouudVsCzen2kAN0JbeBGE7v+roD3usqVWDWlZb9SZFxIHNhXEYdpcPJTyt+B6mTI
/SWkrl8wj5aoVMP3OvauN5vQfs9/kTjayAmSiJYWjXROC1wcsL1VSEs3ggWd6FSP
VzOjP+2/PWHp6ZjAALojse3LfZmPgOg4G3uw95CmXVj2JVAB9tJOVR0CnFLV6o6y
hbU7UT+sSrzMEmADqVRf9igjgOi+ZJ2dPTyN0n0gjFU1W6QhOy4zitZAl0Sj8HSd
Dlc3dUZ4wtp/Usm4p4/4dbm9h10HB0xepFsdZ5Z8NX5fmf1md5ZMP6b3XRvLyyTE
NocDhztqrqcvFjHO1FJcMKsPg7kZT4xNU47YhQ6Ad1z2vDgoSnKIr3lDnIN4RJj9
rPCrlwq46UD6uWzcKbbpwQ4VarXThDdwjS9mPIJbpOQ1ijXN2wDn5BFSyl3zk4Nc
O2I0qRXs4PB3c8RMZ13dkVjAYyHGPiN1R7Qh1uJP7YWcikGuRjFBKgva9TC5yQgv
WnoCsDTtcU65hdlOR/3PxjOChkIy6v5sHFbyL8QFPegK0R06v6EVRVwM/V86UG4T
Ou7MHo25BCPW6AmtM5FIWzxwVF5cfBIdIpMZLoh06SNwTRL5Llg0dwAzQizqPoVV
m5JdPLNtBIwxmaDDViMnesJiO/MKRzwWvdKXG35aTVPk9UR94U/rXTuaKj7Fd5b2
9a7pJIuIHfa/l1cm038XKnq3eTtBPvG5i73e9GwcsLPRED7RktS45EuRFvxzmZek
SkMt57O24yRwNlQ+r2f72nxrFg6mFtZMevY0AKPGik61tsDiH26gYW8+W0Q2Q7YW
c5GVJckKJ/CEKu0njFFQG3nNjdkjKXPPdXUaDjovFPXXrZkxFVwonj5Qt91e0ekf
VzgWtfg8TIUqgewaMv55aI3GGoap0Dz+38RyW1v8RsbR+eLP03SJ2BL9qNcSPWRs
I2pPnjgW30comCEXtZYRsfdDh8Jlfo9svQEWDuApiAAiURqIlQEXDCaaDAOYLFzv
gH39g3x+/bkp8LePR9DSxZnhLaVT4wU9WVc8MtU9lRYimr9gxezk2QyPTPpxm5VZ
EGKKmY07H7GZtk/5/GjgQ9d5J6slTwilfeahhWm1aUpw/tnJw6driZl1l7BG8CEq
uHuYGX3xyv/OlEeWf6SMVrikTQ1111lNn2FQCgilora+IbA2qwLCgtYxZFjRqB5w
80EaOZkc2LZHrFYhteJd8G6Nj8NhXmW2D5bGIWR82Cf4KHXpIlZUDI7WKPPfh+WM
9XqJfXMUpVvDuya4MLAFcRCYt9bYC6fC/oCrTVIKM7TVqr6E56yrochlanI/dME5
eYYORJawWHz6Clwn2Ut0qAMVvVeiPLd4zC6/6vH/UwKiG67CAP3Jwk+/YVZhZkMi
OKyMp9gGFy4r+jyqQRXEBWrjGu8ZtWjEWy/Vmn1Z4aa+rMtLaVHhFLwIxVCfpLB2
4gTBUUao6thyDVe+ylP5V4C8LXOS+Z7F3dgSM4zdN0b9MhE9s8/rGmlYDE89sB6s
3oup0FDmwsrEImFpuKJB6sHwyHDrafNWOArZS+o9PkQeK6LsPgWy0y+6GvI2JVMX
NaqouFDpaOdP5d0aQt16bHktj/YwAJXv97jwXHi9LG3Iwfp2n4ZlM2HEgFgndCZu
qXaJ7/iM+VuUQvFIInhxDuw0FWECF6Ku3WB1udk5Dxo1A7/TL3FWAW8z09HW9c2L
ssgJhsJhj52SfTirF1NaKFZJzGrwPV5BviR2FJM7jSCvNicRTaZsgT/e9AaososL
YAl8vvCWLz+mSMu93jfdkys9C8FHnvKa5g5+10fR9S9OXMxAvSfgGxId2U1tVxZq
OGqROIhMX9Ld6+2iy+YNBTQJDjqirxDMZgka0pm6z5hqMFsJeFaWWIQiFCAVdsVF
JgWl5rMsSPm3iEbEakCkr+FmMNzjtU3nUgwwQxjeaW+BicLjm5h16nGYvQMgS870
j0xxr4zJTWPiIpOkWalfD5K5vZv4y2+0xfyuPdJNqPwtAWTBBkHcN8Vd/mAjR0MS
d5GN34K67m6PuxJK3xvP9/yvla7AtL3V/u0gsh5kxBPkel5aZ5dJ9uTcTNiH4cwU
coYQp+Tdi120aztL41Goj1TGFjFz3tb+CMwj4nlItdXFjFwqOTNUzaDPSH/xLpCo
XCsnFVteW+5e3FV3Uj7kPJh6vW8mNUKC++HjUbDmO3G4FlwDiTcSssP4KoSSs6Cm
mDrrJJJJzylIHL3nkoe/lDd+8abJDDadW/CiCBrGXdQJdpwC6Iewn9c3/W1Xi7un
SUerwWcVSU4S0ujQfzxYeVUxsel62mIJ0AdZI1oigncowIFUTCASGQdqnBjtyVOv
RH5xbMOUTu4K9juNv7+AtqxSa5aho3K4JRP/9+CKbBL6LOhBBz/5cm5jgFtihcSf
EhfUpfzcAqSI1y+hDrZhakg62mwYj+OFeb0YPwcZbd0W+L0S3ygQEjMhWFfimUS2
yODoDAIj7bZ+pGYmYy//QwaateMpGpJnMTxzGTF7B3OcYIE+caUkkaLTNAyrZEpv
PyCZSxhpEGZljY+SDG9d+l14CImbZ+2DZdl9kX7fEWzHDrRKgyoFXHfrvZm8VXSd
XqYjVFXUJ1ZvmkSSBnEnQ9g/YQdtuQotCyW6XgKVGE/5rri8rXtNxlJWylzBkJ8Q
825kIOHOlsGBqVEoHOz6HlQL0Q7+sRYpGbFVnlJdLigUyiZremAL4BObRrngMqCb
Y61XTSRAYMPWijjTaxk51YfBXrA7MwSRE3MCP/OhK8zz8H4vnQ/gZX13c68hc7Bn
Qd2Aykh1E9lk46QSKzJL+s0Q3FVIeqB8f1Ibt+P+YXzQbSRujDIDnXx4rYIHdmVK
cS84UZ3MNrWujrH1iUeaym/hKbCBwr1br+80ArZZ5jlaNWhVjbJpMTtJefqzPEmG
H9zFmm65Izu6A4b3jDo6Wb5vXae6aGDfgzk4RORufe4Ho5AR9nO+jvBVMl7TCZyw
eP83Ju7v+Pfd3R5s4tyA3kGPpPujISmcVz2/FISXdVXGuXGrE/wr7SCMbCe/v7Tb
apdGKOmoZaqYgLPXKn96F2NV998Crj/qyvMRbdxbc9bbEHZMk66o9Z4yht3dJf0q
jNZDH+T17n629VNg4chJJ070n0pGYAzNydVRPBnR5sM0PbgN6knFtI3qJSLEasoG
83fynyRb9z1OOqXCEVA4By2pI2vQl0Aux2zN4u1cgeONghv8RDpH8fVnw1AuFrhx
syjLKRZ83Xnf/zy2GYbbafKOLk+AxZOq3c8Y8tr01riyzrqbCKVdTmOTCgr6+gQY
dWSsBMFFiPbY1RvMDCy6TbNFE2l6HEzlsuYLIh9b79G6c6wU9ch+0Qn11LKdPikZ
f2Plu1ElqsnXWejU+Zg4K/jzhZP2/Znm23yH34ExMVZwYrKRvBi7ITgL9ntcVn1s
BI8ZE0vgCjRas+YpnuXo3C8+MEC3Ik3xCXFJglWy92rBNG33qs+J+oY7P1bxDbxR
1lBlUoHvmeBwSjf//SKp9U8AnCpWRuEfAoqwst1vp4Q9vC88yL5Ft7YzhCw8W34I
vPAlxZr62tIk5bxMe+Yx8Wh8M7omeTVALxCmaz3IkVAwJbuszAQ9QFm27zquX1nL
P0UvI+9HukrugI6HFmyGoL9NN2/6FbSfnsaSWWXL4q7KCpXwnCIc+NnNb9Z10tNc
15bjl6nBLpLd8btV9dScKCL2BI0X5pXx3O16l5vI2viK5J5fTuVmppvXTGQpS6jp
Uxvyq7Q04uusTZ1OHN87X6LpWkJh5gEHEU5Sx1BkIVURvrS2XenuvttyYOPskAvj
PcvRP4ZYzvZhCl+iaZ3IRbRWHJue1Irooo92riOy5+vOibSyHy58oA8szzO3vEIP
FEr94hwkdrNAxevJmVszpx8kmDWGNglDmCQCEPXtdv/C0IZgEtabcv6wWLT7FkQd
AMp8Iv6igs40Z5Qw1hz0LWS3FtUQHu84j9B0Zahxy307ikxPNshB9eWe68W+be8z
t7sWG4J7c04SdMGtzh7f1Vu99ml6or2u19DfjOkpxawLoFDSbouWlI3Re3ZaYnH0
AwzXkz1aPJuzYcWqWSRLY9/cJ8MAIQp6uTRxmSk/4oYPVFIE2g0hj8VmqKbrdffj
avecJtW2UIylb0K40ISrDuewkJNhMNFxDu8RtHrzdRE0ShzSIn1H1SwY3th7SoHM
1Zgmc1M0cCqZkIi028u946o8eTPXN8wTsZdR5QeiHw9BWnAii7S92BWMIL1zHH/Y
5cxWUhbbyS1p2vjzeZr9bNmcfYDVNsmezoiZSjbHcXPP1JcJDsxDPAe1pV1zfUbb
62NfqgzSUiSlqTtqYZO5Bkyz4f/Ox+b2Osn3hx1Wam7/qYewBrpB+WJfeUc6F44n
gJBk0ivaRRdKFSfK4klDA0JD9n75VB8XT15mi1SxDNFdS3p39AYU8oUoCks+V/E0
11PWGMjUzVc0Z5cY72dSeh8d05bTYwVENuPLTBGKuuKSVmkwQqCQWIsY2C2zHDAf
ZuBPH2yzuJ5LytHyBXE3DoqFKyU1yMXGAnmzcb5FK8i4bTLWzDyi/nuGMknbYrIu
Ivp9bZ5TcutHGMdHLhVqOCqhaSsCB71Faepc+1gJpFDoR23LG9NiGaDY92QquA69
vy83w6rULOQ0D0AhyJbWYFshlSVVhaIJuVYbO0Ep34EwFBAIcimccSQ8DVVsZgnn
FWEP/qBR1sUi7mfeh8iI9G8NOaGyIWWGAoslUDhM83fY5iLFHReHIPIEnNg/hT1+
0Cj3L8PIQwxPO78zsZ+GhwQRVE+lZslXKGhY85OkkycG2ufevnh2eozwBRiGnZfc
W5MgiD//7dDwf+NDTzAnxwu6a5li1zAj435pcTCGzcf6S/IhSTmypnv1j0muqW5W
JwyXvB5pgVS8DV1xG+RH6EaJu8XZHkAE9dQzsmVi6n+5KfKUdUZi57pqhJCVCWLd
pvW9JDhLbqE+njT5fRWuEPZGoOmWF9CUSFaR3d4MWsamciBEMF0pOhhEMTYVLd3I
sVhEDRevZ1+5xNjOfjGVdLO/QY8/L0FxO20nN/yY8eE4Ygtsrr8//4Eowoh5DMq5
wyHKWqBQNH32weKACsJmn9gy/3hB1sECIq7e7okmZOJOnEOqAodavSMFUW0s83WC
0jAuo/XRFVCfwSwaLyUgiFRuhyLaGpU/+xSMdM4PwSe7OGjg13pPYO0k9sxGOvJ0
eRrtI7WUqa7hXAOYJ19itJJbPO6H4vTkCaPG9DzoIrFzIlbDDgCJVdDO8pqcFmyF
UTv13U4cAaGw8gtr4JDQHA1Djsb/cHcAyxpL3wE1rXLAq9VvbbzkMy0wU599FCS+
JITQj8pGF94HYnaiozXVNsJT4H77bdNmI2ZzGwWFPxkPEcuqvEVkzmwLSUtzPg7V
xxJYjlkEo8Kgh1kIKOQviFUFMwLv0hW7/uvZLaonN+9FuiITUctHbNpKk+RHtKQi
wZbMZ0DqTONC9ejNKp4o+8Tts5Kj3K+5iCXVoxG1osAckMJpqxp/MnAZBVpqsh8c
EtJtkxnckRPfnFq/m7RclXlP5FASMgIdFHHkEl36EAV0K/R41a0ldQMtoZwq+twi
yFWclwyPyMZo6LasqUTlyMd2N33BdaLxAmnkIEVJl9RW0rJ8rXD7a20b3BC84iH+
Tryn2GcYdwsuP/SA5UuKlNEbjditrShU+qUN1r8gJ5U/U6C9lD70CewFUPi0GEld
RoDMY1+gDozsDnO2+pVAct7geJbuZr+2JaDSpHkt1C94u8ewp0NZWlklvMIwa38s
jKRlKKenbO/cpYarVEyUGh/QHcJJBWTxtOVqarQziyT5WddnQ/qQbc1sqR8wAhtG
U0eWqxgU3AfauBNKZv0Ewot3OcvuhD82urjR7WtDfv43JFg2GIJ+atC85WpwRFRw
pfv1m3rw5SbXDHlWco0TuqTM/5Iz/+XSymgcKIuc2SLscDCXjVudJSXCvNf7Y7hi
aPOQFwNEm718Suj1dZpZQ2euALB6L++/lWBnXAFkI2a/x7mKWuN3nykicpjJe4dI
aKHnJgPm2kOceXJ8WMTlf4qcp6Vqmne3sL9YwQ/ZPCbTCz3wXBEd2xWuJaXgu9Ed
6cXn3AOzxooGpuIvIvMFs+bJh+CgrZnOBL6pvWlOk4OuuWhQtSFQtl8NO8MYeMe4
BCgsTW2UnhaBY2AZ5decJ5mzIUOMvzqxlPNvqyKMLs4i+TPAJ04yWYoopqGzRgFr
koopmmHbVJ+aO41s2gOYTSATw7d+uaapB91FFWGKzW9b2XfdJUQ3AxQ3PnaK1h7s
0grYsxsmBKH99K8WB/e96NW9BVg1twx00CEgxLrYUr/bvNECbIBWjC5CHb8MkmgD
ouXYW5ojQm51brqNAHeWQ+OV42KPD+6Q9tUOhWHpxoPBUqzQqaDZJvjzCRtS+O5x
JEXk8OiXQE98LCIi/iYOCERubJ39lk+Qsj5aX1mWXihYZcfDPralulikc+xcL6GB
5IM+rR9SNfgZl/ndgxf5gltAP4/ltd+noJk0eb8QjyUjcOiDVASnIyRmjaf/1XIG
5nQH52Q6zl3xdZ/4HmZBlpgarR+TreuWNybl39qR6qpyaKXnHda3UVR7uyGRZV4D
f0PJJsJTw2flg7676auroVQ1Wmu/FdpkvSJpgilRpCb+ba80RyoqeDAXFoEJFRE4
PqbGXtDyd/dWUfJJwYxAkPAtCc6QCm+AIa3zqk0JFpaCB2s2gsPlBugh+zxCV02V
mGIaRImQ+W/d3oPOE1lMOnz81FkGzlY0Y1OTvf9Y4vFQ9+fLPsEWughyNsHHRXgS
vfcPg+T9T4Izd6BlIZoHJVswZH0+hugSgkXMmphTPmBkyrZJqi6LO3IevhZAQOqj
NflUhH1B0Jp2XpmfToZUcrWnaVcACinfMboFVIodzRYRpIlj5Qs2gy0QIkvre1qC
ok4wosBAiHxxuv7S2nPIPvGae1ZXgmmJEArMgWaMzdRkFzMqUggc/2oZoeY6a9Jt
2waJtdGwmIq2M8bzzfyrj3VxIRLkIaqBo5q+ahYPHWoh3EvMLw9oKcPZcufHdN3m
/GV6v5JiXLHLHgSK8cxss12Iy2QcJSGYdBsEEEAuyZlr5rtFGeYQHBI9T2CBYK2U
b9+1xXb5NykGkYc9BASgB77dlDO2gV1dyqQzJyB3nDKPBIp4kTcglhiMe/KVadIN
gbW4iKFdOM0oFKSZihTAiPqbIfZBt1OAKLkqcn7ikbcG4ElQKadQKuXL8edasrsD
VjpjGDU72vYTXQ37Ty4erV6NZ4iYI7ARLhmGeCWzSaffzv/vnlglQrSeZXAwV7P5
X+YJgnYD9h07vU/p/qVBSU03LWQ5rOxt2TsZphtBOA/wSoWB3plPo7gIjgqbwqxk
4PeSaqiswnmM3xm8i4V7MPLkFjyBGcfDs+0yzkx0f6R9RjJ40bvgSrITRtDi1ICw
MmJhyTRWxemfqoaWNqG7csOKHi3Ktv3NHWd8HzveX6QzwcwQ13IW9/smppnfsTwN
/ZWxr4ClcnRTS/3w8IynOeWS1jCjS89Ju/0RIG0H9cJmI35dRBpTNMlL3MlCREMc
AS4fw+tk3Rrwaohk/LK1Yxl3M0Y9OCA0XoL3X7spm3pK81UV53V56uPExDUlcZ0c
KjQcDlEBvdV7MuBYgENssgCbeul1dpK3qIFaBhtgc6dmjrjkIIDL9A5Q6HrhTwYj
vU0LNBuAdyhwwSNk4DvZU8LoCCcMZkX038L/OMs6Wxm4oxfSISGjOdJDNPPhH/uW
EsWe9AFegNcy5MlbrLPHkvuFAcF20hwojMa19D6QWWt878k0yHK16Nh07Gt9OSsq
W98lslCJ1YKYX+CaaEwOJ4czqFbf2pFj1oHZHt4keMHu4LgYWIQ9VObGWUB3a7b6
/i1brhfjHh2+pVxGP+OjUrhiiBM7+k9aZEDh0SE5+fj1lIgkFgcaGAnAmzoty3Tn
lX9oML7geTBYp6AV8+RS7is+/QtiN7hVkJbLcttAUJQa1ismIXT7brawzdfxKymg
k4GuFID9VLtQwLd31IGCdMb60fKMtfyy5515B46mK4aE47+OdRDdZzxWV1CtPFFV
6Ji/wv7BMKwmuzqj1cFfzimHYPQH0Zej3P4Et+B4PQ6neJkN6l/kvBPvC1X95oOd
Jf0zP9m776k3GrFU+vOUiwNzSMEt8hEK6KI5zXO6mNR00CqKMiioqolkBE3adM/K
0WtaHsbj2hWOu2sJvfNvntfNKDJNHKSxMNv5a+8MJWa3SkhHXqhZ+KOqGPyzQANd
YoFFItVnhi30IDmmDZIPRHI/vD6O26q5v+y2luvcYZCb4xUwIPUrHz+jMewuiRXu
zqbSZzlr1ikbHIayqrfT2CT+6f+Dn09cGGvfrEBXzuIbp9JRjYv38GnSIczgH+b1
G9trKV1/PlYZ48AtbN96/hYH/uEwOsVg5kim12NlrCsRqfLhEZd5+6GWzPm28rvv
rsF7TytU4YCSgIc+VVDDbEb9MwOQCQ1/fqAmH3eOBGuOEXWPdi9fZdHeumdywfh7
tvk6JQBoQZru8yeyczMQDdcLB9I/iZpoLHuRQLQGnt7wG6fEneWpoL0wQXeHrmcv
qgVSmcPaRV4OsbhAzOrw/vganuvXry2q0iuvvLsGVI6pdk1gJQSMRiRQ2H5Kbn4U
nCrqrUEjVChbhN3hnfoh4xKQaj92ho+Y9tg4tB28jUkdBQFKIVt/fe65Bcj01/o8
JEMVUHEJT6Q3rtwsW7xruBYG096OLFKbqClPVVLn0QCjulXg1sBr25zFezdmOXxI
j/90wa5+kfvRIjH0o2hSdXCtKhxeK774WfizJjwuSmsufLtz+kgTZkzq6Ykmuphu
WjctazR4wXApps3iRmIOTRNYbEd5n5fTzPB3VSY4a2VMsYgb0GGntIH6abTT0jm6
UZeZLihE2UkEsh1tyG9S+J0JL00DFoKa/0SkJNriWkOfmK/iiIwN8rmde/Fp8rTe
d53lR1HNeh4nYtU8YX7YdYFSHDtGai3yjA7hChizyNqklSnG3wJ6epH03sLKN29B
MpNC/5te3jawOWakThRSeFtw4Vs4DNyevTo58y+CamxI3GaDrmkALfj0CUHDhM8x
V+b0FR9U1eu55WcYV7utZxiWLdkgxos5vi1B1enGjXWfv2Da1GdxCpV1RuAPUR8Y
dBXJEQfxHRhld83gvo6YLxAnJe5b+0TY7tdEo3aIeg6YTkiijWxCYVF+RSIzKsGo
v9r2+9QUu+YYSTe724rSdKl6sXla4C1FYgNOu74U+VAtWB9KeEQHQO+axI/Stc4q
xteVDgPCrFUAxu99KI6/TncBg9KXpNuspM5TeQTvOKKeWAOO+DDMUH+0hQIK/h8y
PCgtXWGDsMRXyTcIOGH7CHMygehD6NjI7KiDwAw/MprWWJiumKX3pDFHY/F97XlO
O4zkK71vnf9u3vfj8uyhyJO15ptoIKYQjND9M8PwFrO2wQBkx0w/Z9pl0vZT4hGG
3xPg60R0VxhSwRv5otzNrnS1fPzxpaeunHxP2VFniiNO0+JI7YNFKlou7L+EOIay
Nz1KUld5KNwh3kXHKKj4XGCuwRpyJspKgvtwKpTwWmULxlxEa8XoPVtE4pqauyhN
/YjsySwErbTXIEEhaDfLSHKfBO4KV9ZTgTH0YkatlJrw0sYGN5Etc9EQ8GRxZ9yZ
cYONXFk9qA3t1rxVdPgE9MvIeJ3QauPZBclBSD0zRvunogUxhHrL0TciZPCTyKJi
oLpc3L9rhPcruJ2xPHAoOrp9SLilLJ9k6lg0C1EP8qiHsWezKupMFmNT/Vnt6pdp
TDxILUsPIVws7CWKa2CpP45UPZpJlAnWlUVl0Q86Tv9i2rsEWHAMA2fBFT/CZ3Nq
wVkF64Kw1o2qOmGD0goIqEkY3zsNYBIoObgmsbZ8gWUshWSUdOpFmRppGnucoi6i
mLJ+cke7qTpiinadFkhcMKTnUtoB572DufT2KCqVAMQlTbGlAUzW5bcjBEasu7ZO
/+liq1EqypLKSXcrl4fwraY355a9H4y2fuBlKq3v/07CaCHBzxctCkPM2nPQWlp6
9L9lpdy21dQuLP9pwmxNBpuKMPdPGjXPyV7tFBWA92cQEEblwRdrbTaSGZcuSn5C
oONgmcKn+jnR5mMgVB83wn+2veKw6bgzu5i7/ek4PZE9rSfp3zJSL9E5bgXq5afe
JDNl5yQOH3C9Tmgor/QZA12Maxdc4pi4Y6t/AfGnA+WfX7e9tiNrsjCAIjAK4rkP
JimfecvHDbkbsLDg+6gC/UI8ZgXC1ViQXvUrBh7RcyCOcL3hMmbZYURk8V5GDDMG
mCU0UzXkIfcdmSDFZiSaWsb9LRb6pdFye9NCILfOgUfh+vpvYu8cz1lDwKpE+bC2
Yf/QjxbTLF3M8QRszogqaQgZGk3PjwVnLgNALO5V8xuxaz7CbOlVOXL6uCGxzdA0
t9KoyB4S2AAN6GkYSX8v3vhxrDA/XP0VsFvPflNSkVMi3aUpHDBcA2V6owCffNYP
STa6B36b6+WsS1NNq5NdNEHLs6V56QBArGINxNYTWG3tTps2LmC/7r8Jes5WcBO9
4F6YbAeXbZrdDC8u3qR3GcJgg91Zfh1EjOQzW4Orqj0svVuRSr7ulbwULkpOvPjE
2RGqM8UMPKDkngCK+NCw9ttEevBWqyaPcrFxmcwiFTcRuVnXROxDXCQJ80GHnNU2
SDuKkQm26TCnLQADtVKjzalSBxoOsPMS4Hbk/BZ2a9UsEFhKLwavQi8qYg8WFZ+L
FSvY84ntdQBD9FAlUI/UOn3F2z9lsg95OXOKjnUw/XgeJkn/q1aKJNrbEi/8I69g
3A3QBeBG7GR5RuO7FkulgEwMnDEoTaVTBrAnBNYEPAtKvJxbVEC3crXoFdBepZAD
ewpO5G/HmQjHKJbAhIkZm2LkS39mCzcoLdJ67SGfVUP40/blQAv7dntc/vGp48q5
2H0hLFwHI2ZqA54yfHYj6L22/ipBnMuHVU/Jy0j6moHvx+rvdjua5/E1qsyA8QBh
oxrWnFyF6/T8W3f4H+xui4rMtebv81cmbBbJre+XM0poCKekymOtDR/Zf5ZVKriW
AofuqVHacli4iM++3JswNeJjoBOTex0A6yNuU79X7al+ZWqDieGisdJAz+yxrjQI
WYg/RyyXhzYCQTaQhOgX5phpXg/EsTiINlh22xgYasUQkTLV02QrYaXPwmVDHuqc
Gvl/NXbGQF0xq4FNaqwuIc0Z/IUce5LJFRJGiIaTOCrYfx7q/7DpFNVDGQAbtMie
feJpQg+ocgAQDa3NZPmK+6v4WIsoxKnfDRVmYs2TdY9Xb7T+82S/wNUXdYO0Gb7h
gE9gj7mOccoxfbbuhSEYVjCTmnytEl703TWhqS14u0ZQ2O02NMpGe4m4fmWhaIZ5
pJU+5FVEd1OE+UOrGRTA+7RhO99Gd6fazOIhRCtwjBkyrOcWsxe+kP6IKJUvM0QU
ySC5FgfUosnXlpGdYrj8MMiOU2tb9S+jGRoMHttgY3Y9+qtCrytq10uUjvQ1PLKf
Z+7arOlSAn/ige5NZbbCQzoXR0wYjrF9CKRIriG1j93NS61MpHtnjxRqARZagq46
G4IN+LljEY7cW3VBw1gtV8fvfL8tYr5rDjIsUUOf06Wtj25N9KN2iokiD2STg9oG
6LEKI0uJ4rlLBzWS5IQurSh7iwJHJH/VKfYTOKLnkFSroVvg58n/bp5Xzh8mTcvK
8KHS7tL9jXvfRqYoRUaL7WFF4W/tIGRh/fqvIM1VznA6Zvd5xU7V/qe+28hOx4Qy
ZxYw6lGaqfQIwP9RJ+NpRyqSieg0dDfxFfedpWQk8QdIODc1dAygWWyI8nSKvCY9
3IhxhkdJ+WE/yzQWQlSWi/ztcCaD0rlkNzqgGuNeA4DKpTwdheZqSv3m16tQjPT8
PX+/StuO7+WZN1pr4QUmHtTotMi078yCNGShqbvUSjcJ7EF7TdxXLnY8BBBRuTA8
k27Rr78/5lVqE9oJmXt0hgv2m7v7L2p08q0G6WSHrIBFO9LlRobJ/G7lK4tPqnK6
oUznQ7wLQYoSTeG4IgdhOw0ZAAz4MowQssBLQm1MWH1Xct2Us+mob27nV+GN7Mq4
Y00Gc2ioD86Ll5q05q/rkuedw59+j8VMpKycpst2rymi5Mu/19T1nZnRu+MdWFF0
nJdQbRi45TlCpuoMuK7an0duli93eja1aCGESekRjeCQ0IGWzznhUybMOZq3R72i
9sE2OZxoPXT/UQBDoPoUkfU8q3YJVXgLqYf2FisXMxOGvZ8/QAong8j8BeyVlpyV
osLq6+U8rz67jSGe2jpTdwV4HNxxF7xaqweOOdeNqSm5KkpN83uwmrlHn+K/x2BI
ENcwFeKfpRx3/DRe5ngrmWlpO1rxBt8sXqWD091fJEjCvr4YH5ybm+fqcAM4PvUt
8ISI/f0F2q+11908kQfgkU6jCm77N96oFNAL3vhuGWqVtaYLi98txnIuu8bxqbWK
1ocHkuIih97h5Xr9knl5hWqzCwhGhxY88T95OYY3iE+AnpWKmEjVDvMVwpzrw6e4
9a6IrolWajoLRnGAyUPq9L7tQ+zSBrG1H7Mw15sIQCLaJrFH4D2L9V6vjagJQkp2
h3oGPMRVyrHzeLyvXbk/4q1iJAvoa+IS8BXaK/DUgSC4xrhfLpxzs9bECiAiIL2C
EoGBL2qXbwsN5I99P/OGrCXRWAf5ug0rdGcnQPxPEUL4bDhIQ5hauGBeYPN2W/Ga
5lg1bHgNmhkWoHGCtHPEYIjS5qbYFsPqoI66NEs34PCoOMWcdkgPzEW2kGGbs4I4
p542zIxTKLAS/X+PQ5BIXCjb1ar3/vymZROKIKNwveshpe+PMRmhuw0H6YFhU/ox
oPX0fvv6B29GGvqIhKAAFMF/aZJfUWoItZZBcOl/f5bcLqaS8+Nd5Mhn8+cR7ze3
PqXMJlYgrmsp8TpuG/ykbNYaL0G5kil8t9z4r+ZrpNGjAtHXwYdHm4lr+riRqdsC
jVdT5vPZ2bj712J531+Z240DiMrs0SGFFFv6rnU1hfuPiVWy+FLz6BfvyQi3w9+8
vohDynopRZzt9MbCvELItwl+4HgGbmP5FOny4P1uJ2qqHDARgrFxJj3XYqGSrY8p
GmwMwVj7H5ZibIRXAAZoi/LZHNGduu3bpvbsWmQpM0FlzpTa7XglLIKPVXP3G9il
BIuvYUI9rW5BeNjYtSKJ+grABnCWZI9sQSwBaLRzYexdiDk3jL6uEw30Cp2lodvD
q8T/NpbNXdZKr1KuoqOZLhn3MIhoSycVVTQNrRxoE9FleubRS+YSJmFnP1uLQHOe
mLE/+YCJOj783YxbeBf5nW50XrufmWw9Grz1i0WJyI6FgS5ciXnXXNgiJhkfUmMA
urI5G3xPpWZYm/fmF0LTTO9VSKyLCCXB5O3mud0RN9Mb58fNo0vagkd6N80Szp9z
tUCDX94dy1gGB9saOm8VusVf2Mdtbjkm/Kj6EFHzWMbVeGmVDhMVS9dJmmPPtu72
J5fnkezd9iUhWb11BvS3OrYFuu/2bELEyoFzu5OASdlxigSQTcoz3znfchxzF0gV
2GsURldZ9WYMyfxkt1/ZjOiUyeKWsKiFXyMesOwzLTynhN+6zaFFAUqsxFEOnPBi
5akC1l/Jfl3kUYYxs7O7WXWfWSRx6YuaPlMeygYXMstxMvZdfm8UDFYEliugIF4v
8U7j9J30vvKLFLuoLpAfhdCz+zENjT+vZ9QBIVEp00ywW/0fdGL3VrY0/k6g4B69
4tOv/BD8HHBIZc9SKB5Bkc+ZlYrDgqv69AtDBu7m8sj+oXoA14dXFiSJWmeBkpk7
Chu/Skf+KUuSauU9bVsdfDFikQAJW384XCo+NldEhJ4c83ZHqul/7tmwJRhAKBVI
de4fA77n+HfNZnxI5rzTLYaYcbKUXzntbYuYBp6yIwdJwWARMxhW4+iSRBPpw5ZC
cNwGB18Q4BGDS7P1ZLs4rFBmvxlAqkHHJtSJhmA69Ksxeyaa9c9gTCf+GR37pRGo
yUg/+/ndq8P1xVrPLBCgXWF9whBp3zNLgGnbVtmNPyBl4JhXUy/fbTJ/85EY+kwg
vmFIylFMa95kGxWagXbQkwMOuh9Lg1QAzqiwRJUK0biMlMenxnNbOnhG084tRnbs
ly15M0Y22W4mNOUaJwiek3BDvgTnwgj0OFXHYsZKZpSAkq1XzzDhIJiBKWL0FxiW
VuffNq4V6cDk6I02k8yp0cUSNqCXNqJch3MW/TooCJ7PjUilCp0BpfhkjMHsaHpd
ki1/pyWVTcsr+1Pd9IbQbMf1V+5GNf+CxlZuPY8vy7EgpctOqRzlnJY3IJYubpU6
tBMcrZt+fiD1W2PE2PdJZ2YKuZxvR14Rfq161KTvoxYm6qtHrWu88wgOMTWGlVWu
TsOJlN8s5bKD8H9EUub0vwguRVvVV2b3e6NwMuvf++RBblRzHX0KSJl4zwSR3r3Z
mxFpApemMeppcv1Ya0QO+b0cwVnd3gSGoTtEspfOXJR6RlOYUjMpBnYqKDtYFiW4
HBnQONCAXhTpyg0MD21PcNbfBvtbn+nhvnFlcSKxMrGOFsjFOxvAGZWCJs0XkOwv
wi+nkG0M4eYGvAbXjZ18AKbR7dkAhVfzb2OkXPZjPTQEj2NmdqlNBUAkZFmqVOpx
DTIl9BQsNtZmcNlVtv/5RC48wr5X+6g/BNOcBnUyS6HrfXiZjsjZNOLLGUosH17d
2CMKp921thHB/eWPPFoCfp5MMAkQl4qmZ62+cmxd3glQVIzuHjHS+twK6Xdc53JW
cg8x1a2RKZz6eOBPn24TZ6KMmDAfkTeAqN3ktU+SOEl0cMQVcQyLVfRdKvaQmcDM
8/is7/uw5+WY0JyWY/yjTpvzI6vCZ1EMO+uZSs+8phkobsUdm/p8POnOtQqVLRj1
PhKIerHPgKnaKmrzoh3pcE7MWzEBWub65HfftooxrH2kzqsVyV6xWBx96W0q7eTE
GKtGw/5VZ3qg0nxux21NWDg0AgGUEx9STXguvLB2aeM8fituUntyEUU3xvRHy7RT
QKYFx+UdIW2vyvuHoe2tK1GIY3MU+NwjebqTyK9m3NH0jrCioPXka+IeN9fjKCwR
E8KxBfEW7Rt3qwju36YWN5Z6BmpdnkEZyewNNlJ9runixpPbKzYZvIPCfcCCoEeL
rAKFtfF5gL4uPGpsUlMtSypZF0sVb93nOcIykD8GFBt53KnCDaCvTy8qNfMDEQid
xwaNFJ64/byPZpIQMNlZ/HDRy8WjOPQfs+C1/B3JVW6B9NeUt3IjIBFzBPvzdAEQ
UZcdRezUGBkX79wJa7gvBKIT0YswsTwHAiNofgRhrijPrTE5YI/No/hXGuOOw9t4
cpAWYIG+pbJSYzQyz0Pu5QtyYLvhWFeB7mP0GXIA0hLxW/h5/kVjZqMlfux37qLR
7gk8/Mu/JpJ2ul9L8d4C6Z/ka1yQ244kBu6g+nTbMQvqEYyRkSALHTn4sKFcV6dd
VbIogwjbCZbWhhn0Ef2vR3SR+c72plX8eJbumSYWa12Z5EZhJf27Zi5fClO8vfnG
I6xkVNxKk8H4Lyq/YZmrawcsp3PSOltTO3sVKBrGjWb+SHHvRiHkvdvPlwW/W3WR
ZGMrk6ppebMRKpDam7yzGBTEBb/bl6EonaO+0y7zzmPC+ybCFvyTDvOj0IbIAdnA
KF5lQzqHvogHcIr+L8N3bD7yaMJGz0kg+j9z7eQVYX01VnsT/VfxSz5El8Bje4f8
GkJWrfPaNKtA90z6vZuDaghY/gBHPeeJ0IYXgJDQBfRlSHLlnItge2/KdSN2kbJc
PZzN02hqtPgfEJJVV4mahc2GbDCMEl3LF+SR/IMfe2/3fgmUSfnYWRc0dTSgaCSj
HaicvX51To1Wzwts4qGQW6T0MZuEM4oa5huDzLpWHdY3EvB4AgOtyS1lRXjMraCL
UEIf7g02dXYDoV4bcIMifmKplTDAFagWPeajqbKZ3izdzFCktpzdx2cNO7PyXe5U
bTSzIWT+2qCJTx45yw9GbvjhqLUOS5rrW/XP3ObQqi3YqX5W9mJtjQR8sMovc8Ex
FrmVnJqQZP3+l/xDNZmRYVoGCyjU+ydK7YguXZ/DwObv2XKNs8EqfiOeamToKpjt
fQsBh97mP9q38hMtUcn/gwIqQ6VtoIJi6Lcpfc4/e1mlUbdRxuZWCBr1twlJmkxb
vjO8JzUIy+FMTRR5y5wftJk3WxLMyAz+iKx2cOJGC4OOrGbON1+xC8MAuc38N7ik
iVqabaKJuWQ7z0b1/XAsFl1OBqt3JWdwP2uFoUrUw2UPWhlyGVebOf+SUJep7wON
FVX6dpi4BU3un8MugzFVTHPlbLkREHwKodN0DQGE1XiIdwmId6/z1wwY7Ptnluju
XAFXHOS2YsS0Xez19angsme5CvFMgVrLXDwNjqFKmNNO2X5bSs8AgLZW2M28rUS3
Q5Zw14IQ+EZMZiCTQyzmEQvoCvU3QOtWbV50htkOta5lB6/SYFzpjZUibwJg4WP8
9k7YQzQ8Q1cN4MNquWKGXUwtXOUhp6wtNHDssSX2XWY5OBLn14348gX3TMn5a8Mb
7sq1mvO/O6JhAiH7qpwhxPviFhkRAv3xmroqLiFZXYnQhe0CQUHUjKE3mZhzL+JL
99na8sL5u24PbWqBzHJLuU+KwZSS4XhSCCCI8+4PlHKJMUQYgLqF8Nh08mUn3qtv
gyZm/qiN7pPdAN2z4PqI+kedmmK7RUQCIkNt5ZeuCWz9zsV5fDXiSi7yKdv2Rx2e
XHCGRhh3w9htE7wxZ7ImRQwEoh/yCP/BinEvz14ZEuUSRwu6bn4HMsZV/ucTy4ke
383kyvVCDS0XhYdXi7kW7CI3AWhMdX2lJgoGr7yOOWQda++9HR3+ygFGRuKdd3tG
St8uTLWGwxJMCy/5M8PK/d2s/6DH/hmDa41dcHf5dfpn5Dq1MUBiGrqz2RMPt4KG
W2ZAphtrqOozDRkEAyeh0MX/ZEXcE5qMgI8Xb4U11L0u+QZoDe9HZKzpvw3h9mIt
fLy2yqFejaSpZfWawJhlO9U51OeLxgjnpPDIvzamGpTUaZ/M5pU4XWRmTjd8pzhz
bzfsLHt9/MzFGofySqQ8IbUI9yT1Lthu6fGWAagsAAoUpl/nGqShwo+GKdKDIL0D
I2pBJ0jpZP7HbLqcn4KuSHGVdliR5z67lqQWGPVE+NlRJUb96AJgiDc9JpPhHSZV
FRI+gUtjMdWD0894aiF5quhqZKxWoRdOHmKTFtX1OpkXrZSn+dpTEGB9NuVl7dYQ
cUyAiwMwjCnk9Z4cShaV3eb0I+vFMCoVizwBWDrgB6kH3QNOCmar2gU5rHm/dOoc
XONNMbccWk6oddwZRcOWzQkYmjTIOJQTpj9XExbDJw9jQxmOFea04Nh6CAeIw1e0
qjLQvQfBj2rkZJ05QqX7eKlPEEYKxKfa6BvClFGU9BqfHZTGCve+IuTQmTp0tGPr
o50acTRMJQdlKWdEo/jc7O5klV9ykKHstzZ8n8pb8ZtQMeNx7Jx0xjbn5oGh/GK7
bTANc8azVj0dp6F/VsHTj+bT/M5fNrrcNjFFpxxeRjwTDLQuL6cBbtJUP9jHnICK
381U9xPJSkI874+Ppn7BJh/CQZcmPNV5dY5T6o8UyfQNgGkNr3KWOgJqojSJxABY
GNrlygNi2YRovYuIOX4fAvhjZ0Btv6TxPcL9oLdTqc2eoXqOn//LgLRcv5/W4F/5
WLmet8EP0lDxelNodm9D98VQDIpp35V5fxLODxJ0yKrTIi3Af6+Qn7jxtcdDvOP2
idM2YUqDZTpFX4QOJFQwgWK4dYm1OWRVxml9SOci0Z/sAkaPx2gV7+wCVtHG7DYy
Zf97Te1eClR9QUgKsAPWVtFyRIaN7Vt6rW4C0ILlIqGzNXtMi/YKSXdx7lyvOMNz
QuFQgPv6AHFcSCwLduBCa98fyQ1+3LZ7tyPdzPqJB+KyF/vWspP8PCX/O8GA25qr
Se1+r8OiXzuTuwC1TuklMGpj1Tek1KdFosELTLhuTD/Sm9Hk7lkB/fVsI9TGRlbM
fyFT+uaJqtg3iqhl2YyKjF04X1tQpGpzH+JY0IWSOTTaZ/4gOHL2ufjxm7vZVFoI
h+MZUryeSRTVKq2ZDRahHGWTUot8FP+5qZvB7DeHMogHHtve1fHJuanFDqwF3W1o
gyG2spqBNp4TU68w8YSrEgJkh90jj9DnDsixIObkJBXAcE+bncOIxISUd4pvm++q
hEQRO2++XixAXu4CdCYwxEw8Edrjr3gXMBl1HJQoIJA1GCjP9mP1rTv07+SV5H8l
dqXnvdHZ6upjOSuG8NDi2WfWYnDhdiwSxgZPHeV2tV4nBNOjwiBhJXN0zUYIgv34
gYD3i9N26OvQechT9Ode4RNOmn6aIPLCxK3LGlWiv+YbV5/Vurg82g1F9p3mM7gs
9/jQd8Can1KCksy7rTGQReAq7TxVACYQoSae2+UoObfX4kU5OaN2sb/x0G9nyNZ0
TduydDTqcsl8nkaWWcptj40aMAw2GrQQDQxnNzGj4zgrpk6jBNmO43807dkO33j9
QdR+eOjW8tFgajlaUo7Ugu4csjzi8YqtB+DoMOPES1Mddv6JlIfcX+a/SkrqRe3I
DzGD5akzrT3rv1u6pmJV+hZraivZSRzUYRt+sEDQEJu68T0QUtQUsYXxaXbvLYmj
hcbVc9SZ5/GVka0BeAOpLrhZDKkGXPmFo3eNa/t7N54yG8RDdBqGpp8g94nfrDPK
XehJfP9lgIiAN9v85RllBra7mfQkMTN29dkCdMcO7dicEq6TlcowvJ6sNOV8IG6V
i/qz7XFYVWmgxa/s1Yj2xbioQOxdJk0u88Q3c8UEeOoN89exz2SjbJmyK/yK5Hf6
wexUDXprP+QFcwUWZgNlDZfSMGamaO+b278nsqOC2619Cpk7ao2oa5tt3o3RVoVA
fHkRBlOhNEjKDyCRlIMfjCrpEMhC+v5tIDRXr+HHcJkyopNOK2KFWruZgwaRSy0L
WhgAd9imZr/17ae6cqUg/yWrnGwLoqt20S6g5fvuNFkWVJJ9CadrZgtZgYEa9P1m
MWQtMSvb+O1lv9B0aWSYft3DD/wAXNYkNR7KhU+L+m7OthchUdpf/FXU+Cf9ceeA
1gaxLMR+Ii/FL5+Dp8x23fnn8ihOI2Sp5d+naozR2aIswfBJ5iqEGESzs5AdKP75
S71C/JT3D9aPpF8gnj4GOBNdcqTG2QL9TyT8DF15Tf7S0KwPzKZuo7Zs2R1u7Wm0
dPv6y3BW6GW6XnQ7hIBHx1DMVIajhsAOVY0SBPniWBmXED4NDHSHwYVrn3N+kQo1
PKR5C1iwqRK2guAXc08e9dxOIoQ07Vex+a2dXZdaPF7iwhtGzuGPKGZQRPWik4DI
85+YXZqSxVSkHB1FrSeVGJlqaj5Kh09/Ws3sHgiuNOZ9mr/D0zI6Zj6zH2Xti/xQ
sy1BUlDyganllsHsUIuQ3hSjQ7x5jqp3yP9R70hA6tDP+Am+A5mOopqP+j4LAk1Z
QW6V7xbrxtQlkXBohvrdpy2qni+hbzYX9PykOIj/kb6nyyvjYSlqIhg4t+0a2JW/
WkIuV/gT5SG9QzqUsQEaLKdRoO/MFKJ1OSj/Hb2jzeCL0QGE17lrFR+SkfKwJHSH
pNuPEyjBoXF0MjYItqP4ULHUf0C3NPLLxrbe2/88PLJlC8vL4BUvbbwU7S/1cxY+
9x0sNM0KqCEJoDizQhWTGciVdm4EgRW9citZYpXyifCNn8U8vZKei79gtQOXOoIv
heu2iOR2gHJ1UjjKSdv/Bl39hpW6k3TeQzLFKpSzHGuh4n3zvOu/P/U8lk6aV2nK
tJ1E8hxzarI2qV1V5/91KmuEKVbqql9Tk3uFNgbn4VBV4actJ1SLy9MskvZJvIRy
BLGFXLHIfZHiAFADaXMTUkjIqtN8WHn7+qyG439e8DgHNoBiPTX4ITMktlfAkoKQ
268OV5kVJcHNSX4ga61+O9w2CNvjx8gJ+189oxscXCHkCMyp5Ql+8I5Bp0+meW0J
SEX90OPrrBtUysHb09C0lDEn3IeqgTf0Kf/LJJ35M7uW0niOhmv0KSsAl6EGPGfo
/Xi7nPS7ccrKZTTRJHhVNqiWHj7W3g3UkS7KBgdFtXjdvD3glL5UfxtO5KpqCpPA
zwp6Bn9duu3O11cJBccyyVh4EGfzi0rnSllc+kDDdGotoZ8utTDOf///SfokCFBZ
MQD3Jm4hsWRoVHL0TKXMqSSLSVhWkWct01neZpyrIC+QLfSxt4EAbC58vve4K57r
7T0nJoZxKTLNGZCpI6kB46uAvlHyfeTTJAW1XcR71ODClqgi4FRtLBwNZHBOHAcG
jx+32zLwEqmjl9nIRJBSe5hcJIU6H40sxk8Kz95Ki+Ozvr3E3Db3cf7J1pwmyAis
gerzxsaNUTe2ztjuYz9NdKaiwhyZh3oe9qErNYPvMFNb2k4AnZ1C0CkAmk6Y6z2M
8FxIyGEbGY6vYZI1eFRt/wNdpuj49xV7MCZ+8340Izf9E+QXOH9ngKRk4IQDoCrW
T6rXvUxlIcRSM06MePd/ntSBsuvDv31V973+vprmhushSEistc9tsH6HArpQxtpd
7zAQ0eGXPSjC/0MIsGGU7g37zP++PIT6OnU6joheTfcRgNeHpMcKmEx+Xgg8QHnr
L95ea9tg7t+ShnNH5cbDOtDPaa4kOjO6d704wDb/Pf6VauzjgoMJTF/9QLJD5jPg
seMeF8VMcmOxUO4hWeapdHdNk913yWWdA2wuPX63hYT6CjFpD+lh+eOsW8ErBWAH
A4S7Yuq61zk32f6RUflUCA0jyWeyWvJCKaq6b3CXu3YOx9dx+BA+oe3bXyUA60ME
hu+lmTsWDNhjGcTCg65Wf3yPEh5zIm/OxtamWk8KrrPQ+PwgTsLDAXaZMbC0sQCW
xHdb6lKL/j7yBzH/+ARQa38J+d6zJRzUtj1HWlA0G2P4O5WapoW89slcWhRsDA4E
efhfNXyqwFtoh3aRKci56/pUtHzacLjPBky76OI/ZRkJx1ekl2IJB2ey/4UsnDY+
FhBOcVtIowpJDk6PeJ/Hxd64+AqjOXh+jGkonXVYthSwOV7sk2iuNIPyYnlakSwn
pP39flgkL6XlUM9b3Cz53kLqRW8q0jAvPccdqCuCrHBRBskDAvMU/QMWXA9N06of
dRgIDjtHRT8KtJGg3Fek5c0HShTOt0jquYkE1P60I8dmzssh4eul02mVJhIGdap3
5g2L4leM4rd1N6QpYcYz1yRszcxuReAffBFDfJ2zX8DoATQ0FjH0QNkJyhCSA9aN
NQ1FfOEus+Bv+dv5R9Sp0zo+1lcp9ubet5J957EE6Ew/IAYofjn2q2hJoFsiDc6W
JrCW1kEHPDAHBWOIflPnadVUwhjomi6ZFW5PU6ccUY4eupJjzcdE9NPXi3mGpKlt
j4Vw/M9hHyRHo6xCIa7VU5GVJBTvEsg7H7t1ohNbLjHKKnFOC2kw4+xu3a62U+DY
TQG05wU7qpOTXfZE6D9Qf5rkyRhXfcwfXB6WEOjOO7iqtwiW8zx+y7fjoG2ZOXVu
2cdop+3qeBVdp4wWzaUT/svUgs12nhesaBKJivH8ygKF9xBYZtD5xF5gNJnnbJk9
REG69nyIMjryPvee6A5jCVoz3RqWdxveZqtEY91BLEtQt/2/61+ucnqoS8t5q3BS
N+kbYhIVPCKVR6sWGftwiOBChLvsx3MAmIFgqbsh363k3NjEbTOrzHVYCEMn6u/n
+CQ5mDwjeoHVTp9Fh9dD8QxHLHIOUBoP817rFc2lnnTjgda2s4BUovr9hiXGm1Mr
E5XLAZHVYSiBD5XV5DQ++WuDDYc+cRqCJxqZ8njaR0+b5RcjCmgS4ccSDUJTymjY
qMLBDbdXlMiUdmZLINeAMQHrbRjG/yD+4BrghoeCh2m5ZzJlIZgKSOmGIHnf2/Vy
UU//5QbW2nYkeygOb+ccqVJjkzBzktX0eKGHiCMBABWOEkXo2tsWIw9csnQrl/ls
0RnOg0VdMeke1EzTAgYRIXje2PfP5sizxZz3L9GTpVQLabZFhCY+StL1dsZoQ65e
1A/nRtk1YkJ8vyevzCKkR5LZToBXjLjIyyO4gr6AP1LUWIMxnKaLLoWhV7pFedc5
OHUNjOY2lk96TD/wTWFDZ+YJy9G1mn5V8YFtia23f0ZVCIrNgb5TO9f8+R4dz8z0
fqH8sNhUFHSuZx7a2Kjcjv6rJLZWSQ2OLGp1ry35tUjDMfCs01hq3BTanfMYfw9T
sjgw6rH6PkxHgTygGWrVEaAIVB1FZNkMl1zb6MQeFjAd1liePxdZ0fIo16ohLj9J
ACrw1RVqP1KVKJ6xeB8yOIcr599fXwUC7kNXVmlGw0KqQOxGYlntIRKjqbJTYbhe
FFwXfb7NSYnsfqA5e9k8DA9r8UmnO2kvJnwP+9tPfwq5V+HbSUrpKkw0V1+dyf1j
ps8e9Rgcs1wWumlm65VZzqgXM94lADH5vPEZa0+0DtDraN9UmaSyVMXCSL/j0Q+v
gkbGsJ7ER3dxLwimXDgmAi3cT6kM6ZZnPZddMQqOSaohtBIaHIziISxpR9+558vQ
EtIqVwy6u44UwGPyIx2qissb58iJBKMeGF5u13CCE1ez+ksOJVuLTDfTeLKmFzaz
nRXJPBdcGcvD7Vj7Ka/uC6BWV4fEvLXcmG1DTFhKfePnp0xaTq6xRRFO6QYjbUVQ
kHxpNdCAKTgC8DyaJO2MxhaWgSkPatHtj2E+3zb7uKftt58cst8pvHwBQl38OwGp
Nz4afpQUwYIUblll1sSHbYC7NEMBOFrz3Tl49vmddHNIID8O5tzl4+yI4ZPv3VDY
YopKnxaYsxMhWG9wiHCN0RY6jCTV+IclECcwY9fwy03IempnNPcZFOUoDigmZ2h3
TqtfxSroPByWXYKjGrye4EFrUQTdvn7cRNerBA1HdgiAXPnHIL7fpZDIk9itlRBB
0vgbm+/s71PqboQP2vZP1CKAzk5EHbJGMAwzm7APDuhs52s+75h+9L+eBDXwikUF
8BVHCcJaRHSG+/d8dTgisucll5McFVtvlp45bTGNGJ+rvZhPThECbVbnKO5WQIj9
z/2HLSFL62FhjWWDmUQtfORt0U3acYf3o6uxSdnfi/mv2tK1jRgmv7h4QMFLGTmB
tcXo+kw65WxZCRn5b3SWXQqGP4SUbcH9q8jReiAE4VWEf1joy2LD4j9qeLwbm1ye
ly+g1nI19vz0oHR/Tgwx8TXc02Pd+6mOY+QyCKQX0nTZL4FkckBOD/w3prAikGZ8
oL9wRcOIxakExGE8EonF6OWvGuSx+m2e46BLoxeEY8Ql3N6TADiAQ+HLOqV9bQEH
hjHHebgYSBDF9df3THY/vSOXdOx5BQDXolcA5wiuROVKRaDTrZ3UQEbrWQ1MKmDh
0OLyKkbFUo8cDDdBo1QyD/O0F74YeB+njPfuY0f5N4C0LXjESxRa8xq3UPMYcYuc
VuJKhMkP4dhUqouOfEzhCMFURmLt3oD53H0Z2W+Iw37h3JqFQn/ynnYIr5Znt96x
QEhpXPfuz5W/LOD56W+aJr96OHiCKVVmqba4LNziBYMcyzl+HU+vJtEAldTLLt55
Hod8HhLUzCKOfN+b8vqcfYsyGZZQUfkf08EFMedDfEPhaMxY8fnVfvzqKXaDnqm8
kRsPaw0JvV9HaO8Lp3U1APmnmDvDf2+lz0ZPavTmIueTxT6fFF0iOKBebYxKfhuJ
qz8zF7u1EKoDxbIY8wi6ejg/0lb+uJvGWR1Xtg1pDTL43003TFMJ66myqvmMOyu5
G60Vkvunz3F8F27UooKqSi6MMHylqVkP1PlOk3rbN9cmw3biPRjTvW8hPnKBysfq
lUBop6K9ZnLHtPxMVJ4+x9U/DEEaj/UgAhMVC3aYChF3fgYmaYBUztP5ery2XSN+
Xg2BcRkdezpd9Rcw7BaRBVjxYsAAt5HozScS6Scwm6MgvAuYX6FrdVtvjVqmhhnv
7GYgFNgWyTQVu+Zsx8jd81BTIrmMZP4kDhMuQxWC8kFxyTYn2GXP+i/I24JIWJPM
CVMP14i12/lTlzBZWA4BrgRPe4GOeQW7OipqKmYgNJkJ07yQJIKucPm24MIiRt/h
4knG7g6J/FLUzAo3iY8sg7WbSPsJdSDb6hqs2PwMl6Wz7MDlA6CqW8HnbiUdzagA
Su/+9lnG1nX3zOje6We75MRnR+Gwigi9PFqWx4JG8V/YsmXTwCPUXD/SC4WCTXnm
QFpXVn2GxUBJ2STMrUwv/dmQhckK4dXJauriO2V/vJAa1D3Zg6Lm1WokA/D7nwCz
wckfGSD/E9woOA8n5Isxka/ME3RoPKtYszWUsNXdw9sQiSpnhY/SLAu9T+Q88WvD
z2jLKV+8CpPkwrYgTXRI77vHn0ocHrBJvKZeCBIo981PhWwGZYwGccuyvg4clTJi
C4WBjXsNA+7K2NFaMp9aIOP1j/IyolndSow6pPvcxgS4QbuCQz04QjzPlrlkdAtH
sqM95W4EE/JUFocFdDGSPg0l7mcJfeBZFTDh0WRkW1lxDApqE7FL8BtofmRchyg3
ZFiXX1caAWy98t26LP+znlVlk+mNJadiFJfH5MXb3Xlpu3e8T30/eztVaY/uztjp
KtO8nDbR49LEwYO1xXf26k/2sL4UYoC7+Q/7frj+VcxdqyDsSselW2ICvdAiNvBb
+UdUQdwLcZ1eOQPhtBSHRP0uJZW+ZWIsX9xF0Z7aX+LnKOmi9PYROiNWp7QH8vBa
1MHIX7wtw6e01IBYUK+Pwj1j6J3btMC3EMKA1pExDJkwjTT3iQVmo8CyX0LmSil0
JkkAQ7hKhZYIN7Qabys45G0ulhXSooVTXWhG/iLYrywCPi8kd921opVn+naQnBaB
DKb+/fDfP0xBKN6U8O0IGt8Ejjze/6tTUBFZilZdM5TVimrBpstk2zUhW39Ukz+M
NxV31nxfkEnWt7N7bl+IPPjAf81WEV9WMRXGV67La/YWuSgkxPVzJS2GMzrGcG97
8aLmBtni2EldFv9toMhjLWRxzCNaqhS67MW+Ics1k/9Lq0N6S5coYUSlvQ7+5x3h
0k8bY8wTiIYL5r52NZlfMwYBs4RPfGcvxP7jLZwEmCOdz1sdItzTm1q+gg1bFHIi
c6t38koPRDPNePJ84+rwhA7atYxp/BGeh0fEnMH0gFnqxgkSQYCrY4VrekP5+77d
mhmGkKrWjJ1lXqTFvhZujd0BPz0g1DpAwI5yFU2mI27xgB1SUt1MIdlqmibDHLmq
nZBIbZXQh7HMUODcYNBy65K4BMtgSnOxMnKhCXiqNJk7cA1E9fzKzFLu1IhaDS0W
OXyNtqOHR/jxeCILZE+bj1o3AaEL7td7IZCXaq5sRHAsjXtDNNNYVHRS+L0ppoJf
GSJKlB2vILiCCMbT2t5/9gn0Dh5/jPvKoolGZsig4F/SV2fUiKZItzyux6B1frWG
iPAc3khGVXltRslWgXAem3aTedMQyJx9mO2MPdv2Aj6U/7gJAfQeJqkdBeUeIpJX
V96xG3kjr/MNYSzAHBh4Iohcq4UFDyWECn9rYIpDkCalmMvf8Khunky/+aPo+ATS
M3rC1K9fpXns1vF6dXgFIamm2dyJO9IPZWsnfvFhQ5apteAzRbHB8Iu19AO+u5mt
jLQCYHb/eWGasDBO7WaQkLxfsK5+bmvPe9xansk6CCVM+nel/ZzmKIj23X8V1Qbw
xyaG6lZ/vMHONyr8hYRd3kvjhPoQI9PPNL0nFbH0p6go770CvQTeyVu9NFxDNTqR
tg3T6/e3CYkLmLWXsDf1FdmcGK+QBtBqxnHjbZYQpONhF4YmMSMZyhdkhaNfBMqh
biz+gcVIBuUfCdbHDhQleM67jg5U5wiJPvE9scCLMKidD6S/2AR/Ut2v/tdPQcMX
xPPAM9JSn3s3FzFQ8znb1IKIzr7f9+9ePcfUk2CP4uOMDxpivtG261iNSaA/A2ax
pry41pYIx7+aewN+Is5bzFqGOTwImbeDyv4gVyasLEB0DlMjeq38BODClvuX7hcO
eLcy65T2D8pAWfni0hL93PUbiq2qOoJs6fT7JcTSADb9LVySBFEFVYOEhYHlqHzA
ZppjVLfi74pwlAI5uGKGuReS6bEGddgEb3s1QMFHH8AZfAyOUNLyYba0CeR59Gvb
x9YeOFsjNVzFK8dwwFZGTuDkWQ9GgJYbH/FClRxpzR5CZMixg0dIiFTTsyLaoTfD
kTXn5bPOnxUccAzlqwGyNBufjo/UKz/K0pwwMN3tK0Z3vI+8E27FOTwhuTCfVRNa
mcDrUuMhRTYZBVdkJqvN5xOu4TqnbUf9y2nb06FQNu1N76kPnTJH7fKTB3zEuEY4
AvOmy0HWTWdWs8npBG2nqsLn/pCNksYgv11pd8q7Gxm6hoWCt4XLgbc+27zeT3sc
178GabhKptVgbRbNECOH5pyk7unGvYj7VfqDm54Xd10JgDKrUhYKipFvvtFzrizk
4qZTLaPKERR0TWDMHrYYAs2GOAJcCQjz+MbUvCTObQB8EKXx67O8uabUU11gnffx
ozch0ppTUKDRlUTrdqVrkfUejpWWziixI0kdP3e5ihUo/kuJ7ZysORN82wuo8ESY
PxcICc6XVuPUcsxfn7rMcWHTTdJqzgyFDuMcK9MbgykwmAzs8/TjM1X4qGuLNoFb
c/iom0OFTEd0OcwCrFf3ljRMtas1O5bv4bHs6kHcZQmshejbpEQMxJRJL5dtyKj7
nXfswPhYiN7popCqKwNSKUGvijjSB43G6KIxe0/P2DsL19oeQmGlB2iU4by70JG4
wgL79q2hcdtYe8N2oGkiyEOzizKgEJEaIi+J+o8H0d1PO7UwLv8l7WhOjqms1hxq
JdtoJj1YVCfm/F+dveU14eMcCBd3PnVr6l2aU72sIj+mw9HH0dHgCcqCPlykBZ2w
EbhvdoLSgO8bBVu7LOkKH+oEMIkHldisib38V5SCv1qu9scWUyRyvD9qXJW1xR2x
F/MycRFduh5OHieUX8UYFEFghtB4Hyy7N8kwjreMILtCQu+bFKmdKnWAi7GVfpfR
pUF/TeQzFjncSf7fysMsi7QOySqbtyTivmEMsMQ6VKBNHWpcLLMilqcyH3Hl/bVQ
y+PoBx2ct3zXPQyErwvctNn0pYul4od/oy8Y0hsoH4hWwbRqlCEEUeKeu2wVEcM2
iEspyz9BCaJrZxdseivWNZmtrk1QBwsOU7Vg1+43cre8x16+HoWCTgwofV8QPxFm
X+Oofb/LMEZJNJkUprm1pByndG/P8p1m5D9eoaygsP9bIGPfepwlxAuZAR661t6K
vA4pP3To7e0bNKJYNIoOLVUB0ZgXwuGFSIitDHIPcFTZe8tLx8eN3w94cn6sN/p2
X9cQse2NHVpqCf0QNjaH41xaizYxX17xjg4DR2SESnXy/5HRL0rmZoJpn/KrtaYq
8lSZzzRbeu2Dfz5JzEHARVF4VoTWXFK+cqTTItHmKUtyKqgzhRUjfC+BVdloLOuR
9J/GzcyP5TAQIZ+in3L7bpflH5TiNhRd2uh3OIgQQ/Qy2DnKCjPfrJnSnc/W4w/K
cPW11930blDgjT0I6H9nSusexGRFW+Bic/DPhWaItWyATgo2/YIFCvD6OhOQSCVb
jZMgweJbxVeeFFzzTWDewo+IFKmLj8LhLvrVGDjuI7CLn5ZQrVPWrB8UFHXBmrcp
qGXoy9EPY5mUN2qwaLcBztPL68C8O3ne3m3aE4uaL3qcdJC7kF0azHO/e+hdV/q1
VQR0YVtp+7J4V7eXa2/StG2vPuWEoQ26Yfs4ZxSitorUXSkGbSBhAY79TfSQYWTE
y6XZSZtqADxAVadPyr8yEVKsAreS0w3YzXQEkgmfsclDHR6xpZE8wqJXhocyCgtk
ljSkzoVRhmySAJivMRGHXMc+1QR+kMLwUmzRl7TFa/7g1ao7lHHw009tH8fPP8aE
haI9kICQ+31wSRFPhEhRxvHtf1kpqRZ9hu/P54t9zHaEpTnjMNI0FXUl7Ya8jG/W
MJAQD1Hoz6KJWNnBUvBAdd1VJ8dyR5bWZThFOFUsyOdlOcZMm7fDvMBGlSScJNAm
dX/1czMGt11DbAPwh5aatFfLywc1He2Bqjy6LONkI3NgssBLOKQ8e4FdKchiDz99
zX9rfG+/HsFPhqaMqOw7waHcDVbCVXqSyWLTJtwa5JKTboLjJ/05jxDRUNLi5rT7
XeD4dHKozF4a79KT0IyR/UQo32V/CxiVrRINupvlAM6y1ZnVSbavKqcIFDZK+AWA
39nPOkBpvgdYWrVNC80d/k5+OeST8rEAmkD39eG5ss0d2O7P3ecyi/EzIAQrkRGE
B+VzHpEEJg0cko8gLAAmkFtcNHIAflGz59IRtnr3Vapc3btA+4obgywCYijl6fAv
znIxhMZibPIHmiN/+jZ/2Ip9gB95tepzRdPksvBDZHNEQH6dQ1Zn8GxYa9B+S7El
VPbV2SMFP7cynEJ4jkocJhEuyvv4hH+Ij4Y5Z46KuGMbn2FhP27mG9s3naAviPMk
vQN05hvDIcVF9QWm4IX2TCaeJ4Ad4cXQVgiQqnTeRKuBG2H659EwntJExaZ2Ck13
uJC1wVILpsNAoXZnM0jfSqPJ1FhDCFeluvbSiZewfTlO84Rmi0mNfhVN71+4+b1U
KL2+KI2GXSlJlhTzeUY6fMblkOYl/cXMRfKjyR9Jq0yKXJAHCLaCRjo1rvXd+8Ny
2oBQLxz+fX/j22Tsm+o2/5M9CLuQjfCN47ndDc4/7mGFjZhS9eW6qQ4voDraMriP
8s7oNGlSMOCCDNv1om1AKJlItgD6ON0IWbQ0fvPlluJhGWs85iv+Mv37QyCPpfaZ
JZlwgpZUiAi9HBTTuzk9FW+WyuTi7o4PimXs1TK9nPOTQzzUCNjZpzg+6SMr1Sly
1D53taA/6Rl/ygwnrkS3DgwGY6CjIQ3BvSpo5RRxSXt4hrsBPc5Rqcb2iqt4oAl4
lFQUkNQuHswYRKkkhRL0I6bNYnTRe3UGgym4jHkIbMrKUFXItQpUpoAoz2Vwy7Fu
wUpaxuc3BFFdpaVwYK2G4lc7vPZAICIxqULYKzowihVnmHt9cDYg8lqr6jK0ogVw
aa8U3NrZQWx2J5JJSgmLyknagVCASfxt86lTV0oecyL/X+/hYxToIqHrosqj4e1q
WTvxSi7YPHeqbFJN+c4eic+W4Fq1W2ap2xyrFoka02iWocYwFFSewUi/AxOmKloQ
vELGNVMS+U9s1lusoNvBN+0UrogzpDFxU52BmJYtRTCwFP59Cry4sESqVdUMj8r0
KftGn2CnLtfhca8lqY2n0LfaSZRmYAdh+uNTmJn0nIR3RqaOk8kIha+Hc/izMbad
bLs8eXW1ZG9DqS0Wxs5GkhNrk+hD7WiS5QFaGTJuEDyflL+PzhrQHWmAYLu+Tl2M
HOfxiutrwjdxyvdxNgqJCZ1V7F/mO6tgWV6w7r1bPlU5fR6huXxRffja3tEG/9mc
1taZU4F1FY+GBFqHMgHw0Ke8vHvEo523937HO3OoANbIrlIExRSWxk0uwfuCOLhK
z1fRknvUB767y3/ZsjNyLp1sDRy7dYSmfCchrHqgbsDKvr/ExyqFEJV12UxmSvLa
CsDY4/GEeye3gBUWUda2OBlQgaVqRGhcqGgxLjcJ07fv3V0Vs2rkapy8OK3f/KtC
G6q5rfcyrhSIvmxBfnenWZ2AVdcsAWy+rMBu38+jmhYcHQ4CgG4n8AyqyAaFr6rW
OBrCKHDAe55SKtnqI+8AmFmF52nirTe2RuNuVRCq9D9xmMMwrcZSVn0ie98OdBP8
fKPBeieVcFvx9FzgdJyW2Ztp25Qad9ahs/L/RTrWKmSUIVqWowZaDCQDwPICcMj1
XnEZeHRuqYfms+CNoa+DkL0fvT/6DRWH0MMSx8JYy4SSWOLqg5g/edHbXrunFO4r
uzEMcJbugEgxY9Wp+VX9dyBtXzseRqcCfTeMKPWgqGZWWzgfRon4QPpYmrufbvhg
wE/12PIrueatBECGH+XfFbXXH0rHCuHj0hSZy7ieUmr9K31cFzD17phfaLZr3c3W
he7WkbFRmE8cTg1dG6FpQ30/aCx33SMV1EXEoxiby/HPJBqOqJzR0Yi8FDt/Xp7m
JAFDy8ba6JrnKIW83nYavYW/NAJqyrTavg/OeZ/OmBS7feapAJWW3dyPwDLvzjkJ
pu74U3vTbzEvH6RxENggJen34S6GRQhKGCxaESnu87O+aIDHegWV+07TIO5eybW0
hmQ8S95J1fLZwB6/3uXglelx9MBQNNCKyiuWBgRGJEUptWLBRX1DvkfoNt6+EkrB
Un8WBsiIec6fTf3zq0F9/jYz/IY1siN02qmAZFKQRefzspKz09gt/wwev6G0hNIC
XyPXgh3EFYoyqQ0YmfXI5BhZJkx5OoP2z3Zbjgh1DBmM/qhxTvR5bQlSqEti2OPV
9vbwl2EO9M90Ihz39WKbL6W7G8L4MYIreXNIfgY0s9cAYwvldobBD0BGXqctd06M
Bfymo1py+XUuBVqIU414qMSX99xOTg/32XjjBpabiDUvN3ZDLYoM0CXug0IAGXBD
OAH3csdOeM9td3/GlLaOcD004NGEvTyjGeFwHMhfzTxLacq7oxbehB453ywe+1d7
eGN5d/C82erabFjRKTb1Qx0Amp0cmzpANk87b9dx83Zu0nYmH/NaFSW3ooRG2/UU
9avmSY9vJyyXkaldzapYli5V9oMFlPOooJW/HgyxNErEbXpbPq4G41PlhBAzqZd5
xlOFJw87hwNUv9gXKLwrtWjJFBDGznt2m1Gs8XDmY8DdGRcXonDYDBjtxEO1PZUG
qFoEWh43JAmDq2hEDPatrqOCBbULy+Dtblnu11CRXCeG7/9daDmHfKIvINfFARnA
nMpJyU4Gyg1gEiWVScfU6mCp/LZWqwR3vKRWq9kEWUxMnjtS2Xsf/+RrYFxDVdMb
RrLm9P7/rB0u0vTT+IvDv+z2I+bzX1LIaOiMyxQyhuAtF9Dvo0IDXvUnsp+1opE4
01qOO9uQ34NNjSJ5KRYviUVy/5BDrmRrfMC6mTzZUS0yNHig47IVZ+Oog+YdbJVA
Uz6ksFLszGN1YkcDDgqO2xqcy7nju4swmKNBdZkvu635m4U0WvaI1UsOABKhOpDj
l3qrXeb16KU0p0VdJD3SrJVkR8ICUpaNjBDFCITR/bVo3YhDGAbo9/SJYg3I1XFs
DwdgcR/V+8y1RCd/38cQabL2I6vUlLIyhuvf2VnN4zaNX7cS0J4CHtr/sjN/C27g
R3ljpooZBqbNF+mINUE09SjJQLjr98fWosEfK8Tc5aLtA+LuqzPq2EOm3gWgzu4T
8CHfq8RfIZynGBNW/f2R/TBtEfu+Ep41zASg4ypmf96QyqrtfURvBS1GgzUlQ/7D
QbrxvXxDpmb4umA5WnLy46fxoEeTzMgMLTcwmd9/IL1ywdIm4FtTPeOV6QJs6p5w
b3wq+jS1Qa9uel6xzk5j5F74nEN8CAdnjTtilW30mYdjvnt3jxEF2UtpHuPZcYhW
zfvYqwmVP4JZPRdB6ChS25IhVKW+Df2Ky99GuUTF0Ae79CYgZUc4UVufWfUBi8ut
ygojyc2aD/HqGE6tbU2gF72UChMth+/F3+IjLLiW8il9RILeb6viLRw/lnHF40od
JjsAFAkg9+XhrsQdtvX8SbAH5n0zW/pq/pA0Frde2Vg4DPrNLvEl+0T2CXuY9j0C
gb/cFSliKRIMqx8W9zDL/EEc2+rSeaWXGbX0lLb8gaCSpz1idsWRNXIeaYf0OPdi
AE6qxEWk3kW5N7YPlX0O3oFZCE6JuKU9Na75ql5V6RXLsJB9i1Wvud2j0apJDr43
TZa2V18H++w6uBgKgARjDn7tVlm8TL4+/FKPfet3Q+KsXLK0bSAYqofjkmR6edaj
hid+1+dysn/gVww35sn26zirY4SkhIdss3dkbLHf8tVWUTW63saU9aqdvzKcQSOc
JSiIT6R3fxGjGi0xmr5BUuVM3GsT7neORu1MM998boIXO0Y4VpKXxM0DRfkyfeoF
E+JxxLLJOsYMkKdtZ7/IJdI62GSa1SmO2zmug3WCCL6iulDrkH5tyK377SOc/JO2
UpfnC0M6jizv70PioCtnivu2uO3eTHW23mvvCVs8d5sZ5BCnm7/V2Nz//Z+H3M11
9AesRhAkG9x8qpYnmDY6pfG6UkRHF9vRdho6LZQdwuoRpEYjgU5GTfh2IRJyJcFU
xo8LxMXw9ovdBCPn2aqgJT3U08Z8oDLmrKwcyBIFQNRZhytQdyOG4bZ016/HQNIe
efKLMsKHoWKtpggCFm5eR4Ukvfez4VCY/6cHjAnDTWnNf58dBHSipYKB502zAeQw
k/uUhioZcgxntpNSsZbDcP06v5rbm32z4NgajvZfDrE+Un9E6x8/CXbFGGYzmtYk
8XY2z6BQ6LbWGGj39gz478Pm1TrVhsETSAW6V8FaxR3SGyorFJ+ThPiRqHppBxsh
qsDlA/A1d1CWwLzWjDvxej1aT9U905AdOsDm+8Bkmc0lSuwaS62bFvuH+ci08JnU
E4f2Qh6JPUE8OexkR/S6zB9r3vj/sigVkAkhySwbYtDKss4VBY78dXJrWnbKiBQ0
NAzyLfOk7bgxYQHq6FewvillaMdkDZPJ1B+SUm7RD+/upv45S1v9VeF1vYOdHo8L
tr2E+VmuZ0uehN+FmoGGNvb4YLPzzZkeWxMG2khfjLfG79Hjw+jTEb4Z9JrGU6kO
ZSo1RQ4NoaaxtsBBmbDmc3shaRoiWDfYFi1dvb7POsM4R0uQr31ugKOuZaKcaggQ
NImGaoEKrcbyGrKmhAbUSUVXZZFu4grXTKxhrz5hV7AQBF4G5sDTZ+VfInhp4KDD
/6v2BqDmG9LTSJqskSgPhbmleTkJwB4kfHtDlb9ja5twRh576GjZOZ4h9zsGh77u
UJGDnFL53Vp57Gfk7gIXQleQYzwdo0h1/gljK+/7OIo29GukujvRNNZ2m4mrqazv
DfMN3xVSDd3+utaYbTzpnC9dOnWsUNIYSvr09mvPrMTdV06VIbrDVCJcl/rYwbAV
lAhOGoY0JbNcGBm2/4yfWUPaCkCyszriBQKkhTtfMt9TRXLHnvkR4OqxuE94mpWS
vzuo9EJD22rkpkPlRmgOHAI+sG9AlOvrWMtPOJWM7SL2mYxUTrNdBPqNlvYqkH9T
lErtABdxVCxayg6PVQISMGk62UcXFae3E5+UHspJfwIgOZPX+Jx8I+oGrBQtB6mG
BOEQ+6LKZ1FFZBenoVHxepy16r9GdOoQ3/uPuO1kqe7Ny9hdEskzQSzwIOWm1NoM
1P4PUJwO85UK+B78EdzR0CT8RWIpTP0tmFfwFdlA1YQ/o6qpCFystO9tntJxVJgQ
GnvMWxIX0sGLn0dLXBXm+MKunrlIrZLFQt6rHaYGP13XVjoOKRDefmAUaLNjcSa+
NOo6C80vT1h0grrOZPa/HxsqFvoGs+TQPziHl7TumqHIBoynHRthNkDR1tCF/SkY
YtcGONr/nQMGP+bKffC9olK7WdglG6RfXbTzjx22oxQeXV8z5KvGIPZCEllDtZhK
0g6zPXFYNmo1dnLaRh6j9qfIM2Dfdc9W3QO51143ojAJPxWw5JvZepwLNtZxVjES
rW6Eogn9PLif6MOD5LGTVsTR0e6IMJixhnbU1hfGfw08tZ/Zyc8zUiVQi+s8wa/E
A3K8VLGbmgjpTS4Ge/7pWLznrD2FAqfTvFWEYWj0oHmVMiQAkLJfKGGGTPqEdL+g
aKWAqNjgp4gA0SxmvlF/Mji8z2kp2OVgMBAqKdkUSnfDbtPy7La15ym/s2/w9Oxo
0OyIzX00WAx1CWJtXbmkr2TJUn/avhbYgEJo07fMJgJimYxtHq5jt0xiVL+F13Gh
bG7Zc60zqzcNbLotuCr7QVOBoKsl4TummGpW/m4zyfCIzL2foDOF/Zp6pfwBGu4X
bKbF+XImeDTHDgR+4N0vBYXDc45M2A7WxiBgudX9o3wBWkz3jsaFOe9DRE4s9wzv
ZGcdmXybsWAm67xXKhdH2D2BE2Dt+LaOMAMrnxQOt+RryCIs9XdE8sDUbeFd1zIX
yZxUjyCYUzImWc9RVPDzugZP06kbdsVT6hMElqBP68jhNsjjy60+qZD+NOsFfZr9
sJbudCv0HHuc2njOfr1ILUcapjqxSbpyvfQ5DvsNxE79ZlqxvpWBu6PXBEHNUhTr
9foTmmVr/a7HbEk2l+aOga+f69BdU03yn8NrETbexfN0+L9l/uCfrRaJY4sG5Bud
AnAyUASVTHHOUR+GB+XdjWXzikCfp/aRhC2g8GPnGqZAy4+Sdm4/nmKxEj+9SfHF
x1J9YK3VlV366yNSX5FUhHABDffGnU//3wQkRTxOgG2MupCG3m5ofTGM+dWyvTpr
1Gtemiu11KJyMTfaRyOAdzDroj9yDJZBmsENLS/QPRN8maA+BeLu8MvE59SpuvxC
p5pNqB1yw+n1ZaeLcvl8FHqX8BnILTVoJ82qHiGiKCZgtBi3HCQnFI0YQ0nKInTL
tEetPIND8n2MtH+40I8QzY37WWvW39uU4WaTQxEBgMgPlcBGbhuOvoKgwQO7jwSJ
Lq/GegEWnse3ZVw4cuh7B7oXFhmeWpgSaY6+ks+LIlKB+iTBhAeJDVp5HH/tbMyE
K4BK6HB2ruZIulPDSFWEvz1xJ8H7QSsdf1rP+6QTQwxJmVCKvIW8B6i+wYEq8Yn4
xRCqJ99nfTEdStWCXlSXYwv/3vfDZDJFn7Dn898RuYHgoMGBL05lBvSGAn6tnqaU
oIkaMo7PokVx7Z68+Y9X92qZKv3QH6MGWLehnNhtwbBFNV9GhTYRjwE3vX3N6BmS
nMP1waqD5k5cK8FnIDl+mWVI2WbNCOR7xOiel5ZhJDDSfAaZrqa35moAB8WZzgbY
wxr43klzTIAUS1UuIDpWiG+SGrvGwBAVyno9eoZq50mf9pDMIDp6WjXkyu2FlAY+
HfZh3crbzCcO99BPZMDQY93oM7Xx4bslzlKZ852UpPnFC1l+gbChoo+rO3CzwUly
3WybVx7kL/hy7GPBh13ZSTzCJvO0BX8I7mlgteY0RDHCUDogiRSzQhs00AkQYjVC
GQz3jJX8HoAw5r0Vx6Njd8IK930oJhcgAjoSjH9oL1dMiQ0MDXC+aMoFJRaK1iLc
ufQhLli6lGDXHyO6chJIu90mBuTAWd2WWy2MLXObunH4kn9HySWhCEi2jq8gWHml
STy5djMcM95ZcsS7cTHKKHxmONKVr2YSf4dyaXvPX/Xja5nTy5irWWH8/d5cGJ3w
SIS2KM4xrtvZlZVQZHyiR5Icn8+E92STEAXAazv31hsz/ruAE47F8PIolxxa547e
3Ce4YtolrDL6ydfogmqu7it6q1vwjz3FxKTToYpuYRL6hEx7bZvTy9DRS4fh6/eU
isiJ1bjQ2iKuFXCuRzsmNWG+Upy+dEOzia+OdZTo0bhNO5VKAK1nRk34bnBG/6AH
SBYWCD3U37mg2nJvllpH9TS4BhYwpOq/qP03TCNztidi3vD9lNmQHO1vBE8Ep7xI
rt7ZCA6aUz542/qLTl2z8jIwnE9xhfOSTzSxbgwWese5j8UueNv6oIorc6LIwA98
ZHEPHjA/3plWq79LWimgypq67IclfbOccY7X6GWZXqpdezedRfZo/FMAEbbNR/p0
aNqYskhs5aCydVgJF+c4ZeHn1ACRF3ke9Cxs0pKjb98nt/mFeHVjcCNE/bQCGDUN
jFAAL3qPxj9jo23OLZXnBn3RM8verKOQJg9OcPYkKhQX64Zud/IZFuuxoZ29ik4A
t/dtFHAhl+v471peqhVeEZ5BkOS4gURtwuFWohWVM0atj/s0F+KpMjen2nKt5XMF
35tORliwHScQOzYjrv6rX2GUAxdiiH9+rW/kcxBmRJeZ3/m7shZ34geWfiamGGXd
mpiFpTgxrnKCfIu/x16+wNUb8Zs3g5nmQcq8EZz4eQOKh4A2CfRoLWUl/xkqvBCQ
HKHhEZBnukQ971oUJdFecEgX9cJd9Y1KUmOe7D7RlwuTQ2z4idEIf/fB6dh6rckV
oZ06jcGZqsMqCa7aOflnUPmxFY1pQgip5QUH62/Ozkwm8t/uU/1f6xOfYVjQLlTL
UAKslN0USyOycaur9sqKP9p9ImZGF4Yuprikxxewct6NhVsf4encvGQiV9Dpt7z4
NHlpVwOWRjCZqj7FUo4NW6ONKJQic2fcEO9CCYI714SQuqVPNA6yT7Ja5BdRt2b1
ldVm+8+/yBCJURuSVnwDC7tmrUg8lHNTTUwGHF5eJVctTylKzRZmx200wcCrgC01
C3deBowK6KUDm0SiMAhNL0jhNZWia9Ga0VrUiwWR5dkizcObDLoyMrP7ZAYFSHCj
XiWC0lWIfeH912ebQVslXxV6vMSMagTi3YXPrpIRK+sy8cM25HmPpheH7JPnfEyw
5sqsuJ7L6USWJHsG2+BtQg8giqwWVk1UQwJ7dxD4XmujSx2hfnKDvq1LfE285mDs
lfU7C9je/cE3Xeh7K4VKxvH4f5apFC/9Pp7IH7Ok0PbteIZcBOzVUnmBKhk+Ir9Y
9dInpUpo1JWooB0kCPJ3AoNZpJxrDwKDwCZugMosQzaWoT5Y5gGMtlRC9KZ5tbzC
5tt+C1XBPmNxTABwweEn1sahHHWKVlETHhdXKfGIAJKAIVlGbdVlNIAbP169E8lv
4dOI3ZAR4FPdmFe9PISLrXb3NjFg9brw5jzvSubK9THyJ9IvuShaYBPt1Qe2oYLq
NjYvFrEoAvA1/zIiT/1HM75aDEdQKqTtwgpBNgRERT4bEEwCvmLznmzyydSYMkaK
ALlHwfGgYjQRjArQ6wpxQIKTnRXbDgNgLgutVY1bGtwSTlo6EPOytWip7cyD45dI
QGxrFelQX6PQbHGwRResOuU9Cw5QU/rRnURSaK8na8I6NAJOOvStskXRpbTrWjiN
4A/6SS6nUE0uCeJo4S5If9DyjY6K0SMT3IkFxQFyrXl9NTVdsJCMCpTsdd7IQ3DJ
R4+SawJ9g7HJhUb3YiqNGja5WL/O2CXOY0j6Pghosb+il8EGxJFRUEfw1TEHOPmE
1qfezRIlOTHbCIWs8xNVFsgNy42Lg0RBHXieMbpVxc2+qGJJgAv0S0dq3N5bW7eB
YROR64nNnC/P1B2gmSzxfu3XJ1ql6hzJh8d1qfqrqDQfwZWUj/xWlcQgSF+Z51NH
31D5krOp01yxQ/mZvnVoIf7MDgvVLiIA3YNBivq/2l/07gfoZ+q78sS5h3VH+Rx6
ut0mIi+b/emztmFrQu55UnWFE8jEJndC3la7VkfuKhM+8dGv2RfnLhYRDMC8sKzJ
V5BpqzWbWPr8zN/U55/Pk19GRY3pHEvVDEl+aqejeS8VkhFBJb62EsdTWwIn8SFo
ZvFA5auNATwE+U0WhR4p8jNBzZ+5B+cJqN9EE+Sz4nb/0xBJj+TD54V+N9qipJPh
BbnBsmnfJmNcoJxAB9hjmPfGIlszdiFC/f7OgAiyqSwSuPE6BLr8tdFb+JsBGm6+
hf3I4tffK3GP9SBCdDWyNYfRcWoWhkCA/yK7gzRkXbBnWRcvRxViI5RVusRo6f0m
ETu1t6hLFiVb2DCn0Mr1OgWqO1OzvG7OhOZW3kp02IYUXgSFaHqmG6JXZT+ZAiWS
fpQRukpaxeQWaHwd6vYQGs2+HAvd8MGTA36a51Wmi+pCYVlbVe9MDf7BNvx8Y7QT
IS4xiyJIiPM/xAHEXVYt/8Zs5nNcYE+Ajk5zeAqbrrj2F4K8fHTcYzfq1gXnHsfD
8A/Lz1+kRcIiUfmDLquvw6u70VIgy14rw8Gx6kHFm/r/hUf5bsyd6DPzqcAACJj6
OWcc8B7ppGV1Qcz/0lR+xTVPn6L1UpQxCCiWcq5zorVtlKcnCs5E/OCstc2lwX8x
i7oydM9Am3sKM/ewrNVu96DsEiJEEK3X2QY8zAczFwB8OPnNlOab4UvHMrdtwTzE
XoeISsCbEyMKcsvLhkrIh9KU0azWemp9pA+hp/+277L7mIrDvFBvUrYzThKBPQhG
M0OoQkHfCQJ09Guc3/KjaF2811ZVd5bmQwsNn30W5HRffozNCxYxXwNROk8ILzRF
ya9C7l8s+/b7HbtpJZlqYEi5TZOMK7smFu7BvcSoZZ5mJmjrPY4HUbsu8kiLqvTT
lbqEzqEy2xTnbuWEzn8GY2wdBj7AchUpQw9UBE8tOTj87zmEVR5DiDvUtg2QTkCU
I5/DWnv889EDZQiw3x3K+X+sbi0rdNnx2WJDyTSDg5XuTxM+fGX2dMQDLxqqotEa
XIwPXFtMLrExVs1avBZZWcY9gDAssnrLKBJSatJmZUgVabpyM6kCvChMbLj+p1Rn
gJP9eqhAYUUOi13SLWLf9TVIJjWlaocyaSSnBOtNdKTOI/AD2DXh3EUFPnG8Th4X
sJ2Hu8GA72r4MyWrCXwwCv2Lfkal3R6AKdtqLLM8+HhQ0S0j+YAlv4hnAHiXoX4S
SwLk1u+WOEtiVSsWMkaMw3UDzr4kXa83xx/kfQG/QA7e42XZtkJEBmi90ewENfzY
xolrPEq3cDIxeP9FdT220RqDlYT0bkVyqkqui9WTQhxi0D5uVejzIz6dNhOm7ZqP
z6W1Bbm7GSBYPrirIotWQtntgqYPAbXfSfI2yxNk9uGnPNGbdRczCY38kQyurO6e
wvgeodPjDxYxkW7H4kP+0TLJ6pguHYoceHryAxe744Gohh6n7PeWWjGRukaV2mih
VHOhcMBV5hI/cFQeiKq0n1Vk25DCRYCWlGZbSs9geVb8q+lYHrssDp+Iw5bu0GWU
fA/CoMO6uQ1g8qwJjdqbh7Xqcu4Rtpq3de9Wu6y4iDDqHT+KmySGsv4KHcqaEk08
8aTizKUV/keQuIHxjC74PMMgvdeD9vA3SitrLFKcOJ1k3Z9CefBLNdYY38zXI7uq
5hgG92l+ToBzywQqQyW/j4CoTqhNJatEWcXM7mNle8FaCW8bwd70H9tK5JgT3H7+
ZuBm8tYOOuNLiVm/PL2OnP3oVwqpvUGEPofBfrK4eLUGVavZa4YNU8PuaH0BNLFm
QIWwg5E4pUidcU6wKOezFGyMiHnNqzYuEsITlOkc/H1aW7N0B+hXjB+tsGeKUjbu
3JW92ww+YbkbkXOcxjd+DXixzcPLg1lvfWI917BSCL+C+QUvZXP1dZvZbdOzaFly
iJufcImFhVRhAGoB35Iu9B3gUcQgLm7KVKBt0q3tpq1Z9VU0b2FDxmWakL7OohfZ
W/EZgw8HbjhuCc+d3KK3ibW/Ia56W9kJd/s6p/0jKcq95aT/CWrG/L8mhfsWEIf0
nw0hEEnqsE2t0YPmotv+yVPgBJGFdfW87J+Oj7C7iXHHvygWBtzFufUyJO3Nw+/U
zQqoM7PtjZntTIW587Af2iWzBsZvH3G0k7t92cAZiGSnbv3uL7d1CblSud+tqGoc
6vjIfD2FPAZ6m6a27rLOt7elG7hJFLHy4SlyWz1pf/ZnXU5f0edxIaqsW2Xo3b3X
1uU8rWCuzxJT6MAaGs30wodgOyz2mF2gEVJBWQ7KI0qw+OTVK4hhRyWmeRN4XUq5
Wjfp1AcXzkIz0IN07AKlGyV3SeoEAo2wlzNjQ6kal2qwKB2KJthKIAMAD86HwLr8
VO5vL8KcTo+LpO3yR/Q9ZCB2Y/ra0EHJZXFZL0ZlFFUCZq1kifFe77kwX+r2a5lP
ULyILX3d/HVAOjB2i9guniKU80T2bNz7NMQov81la5r5rLbrR0nLyqLsxI17MlUQ
TdH5lcfzrTqXGOSTkSw6GDUBWVdETC8WprkneiNJTY7JEm7mbxUCkstgi/Fk33dG
jj6YLkgRpMd8bsb8bg7TKD1rqMPiQoBwlDQxuZFQiawHPveCCvvYUyuentLP1jC1
F1AHOUS7PXHaBA1KQWnhD8go5qd/XDrchjCrN1XOAJ97BYMlRU0ReO3qUb/4hzsR
YpDAdYCtCNchLQ1SAaJ9fveDP6wO87a6bdP9b2zRQIdvxXA8LDktt4W0G0aE/hGb
a89vCa5DryMeBdxx0FbHLSc5gs526k/jDlZ4DkMPuSJNciiCEiiVLJ2vNQprIMxX
UTH/NimiVNb4z6G9w/fhuzmHHIlQFsfbO1yrM0tJ8Q93AfwrbGxU+yBSUo3KcWJ4
v2od+SRky1T9IFf3vzoc80gjH2C5HwVGQs9wkrnGwSlPqsJAiK9QBlGvOl/JK/V0
qDL00RHbL2BN3c/3nBY1nAVhZIU2TxiI4pUJzwHXT1gsqLe4OfwJPPn3bNzbEkTv
sZ4FP5VAjVn3BurOwsxvntrGHS0p+q4KycHSIINNxDZk9fCSvW9EhWw2R8V6Xzza
YkkPDsF4RgqZpUE1kEDCiE9H2ryLp/W++RHQBvXbZa8QRuLGobRVQRyVPTtJKXs0
RdcPIVA091d/Jc/hdxaL/1zIkPfR6SRhVlGdYUq34ddk6jfj1VEphvpdOlI7ZiYG
eFkqF9xJJqht2IgDL+nJyTwaQcskzVXMKGSTDuQCKjxnPevBHFDsn4UH0wbHbd3G
6gdVa6Rcl6+HB1G+iEBPZKDKkiS3koGfEYjNMm7e9eWQ76kBynzGHpLpeuv4WqAB
EtNC9SUtanpSQsWitnTn6M7dK9J1+WRNGwSDxh0jHvSLLSACJ1HZ19O0E+py1RYu
5cGkCR47izB0MVS3VeprctbqtQK48AB3X/dqdo6py5wWmCMrMK3aY+JzPzAAx3Yi
wmiic8PEcFToODlBcRvBFpx4Lzh+YXqGY8ROufZ6yAkHWBBw+f7iB3YY/E1ihHKl
unLrko6QAn1lKMwUKg5xA2dbjhsYaLB8B05+yw1v6G4O/fZptaPPerAFPLR4bgkv
aM/UK/WFD5nFNSbOZZifx3sRSYttNIpV/cG21+9Mui5J+rXBpod0OGCyoV2ylVtC
HYDd9YmCsljhILnXMERJF6f0QMxvzhV/6D/XAQFGlXWtnOwtkS6kl2Uv2qjg9zcT
0z3GouFwvKKBFQll5lLLw9meBtxzZjBqz5CvcrLFDCyP69rA9a8Hd2FG1fYpLemB
t9FB7boqLQuYRLU4cphMU8+G5m36CtQNTUN315mdS5JN1V/yKcpIkWLOKFi5T1IV
5cjQvwRvkhoswep/43jDM1CL9+lkoFXhi2yr3A1pk1t/Pj5EpAyqF3LLbfh3xgos
7IaJdUx3qgFaOJJHThb4twnhloLYCWhlF5u89szV5vjG87/dqWIm1hjxYHcu/mp6
1JrFyRnrD1yc/QpsgeOECjhAEmUJKiorGGERZ2mGVNOHLgDq1xC1YAQmjstwSBgU
JWh6swl+QVm4d+xxIF5KAtvYigwFV6NrMXCKjFZoFHxKTEgLGn4uX1P7HWXkz3TU
J+TRm3DIPYIJShX0YR1U6DD7RRk+Q/wExmCnf0ruuaYRV1uhNckP7q+eBv90VMOF
26knG0Q2C042RpFI525ekA8dnCfZgxB4jlZD9uDRdYP9CGAgdBHKaDaa4MPgjwZy
zcmdcW6fMv4e8Yr+lf1bPBC0+ArxmTobv311pyPGhp8MsX9G88SQh9hxui2kQ8EM
3CxuEIPYZwNun3d3Lx1FP90ZYqU6q/gh7Cap9e8b1pDwRU0DJOrBL1tvDwo/CbRW
ytDBEeDxIRq8FRtcn3vCMPrDbioRVnqe++33GmGK0Mt2PMsw4eJETGZMpxMS9AL2
LKLWX40I7tqiKy0ZUckjjDPzvUa3unqZy3gc/DNdcYnPSa3vQMbvPYvD8lYc+Uw+
mkzRjo3FYGrOefs0oKy0pYQLh6j7ApN8Tr/51uAakcjHRyXU8545d5o/mj/fUMZR
4oLjOZSWwhL7NZ7YiIXyaeOqeJXG2iAdjHvcUWI3Fjf9VUx4udNdKLWXTTMoa/F2
jN5Lns0OEhX8zCfXCpFqZfzblFJWIxSNmGxfpWjoIHz1cnp1tLXemBJulElGMK2c
S5TEBPQNya/tnXWrETQ4UT8ZcYR10R57sDV5x4rtf8bCpqLMxRnE8Esg5REbHZyn
0sfU2m0WP4yfMrOGNfAVAlVzUSkA7dZaAyA9Lq8Io/B0YsPIqD4mdaYVX9uK0AVp
gmEsxQ3R9s2jKOw1WbRtAmbjjjqXJ7pjjJ/qN6FiEFwaQGXyVOW/CsFpJU4BKfmW
qKGGXxmj1T50H9bualJosll/vMAzWg8wx5Nqxnfrm1Ckn91ZlabtmZbsVYwYPAVy
fqGjsf47xci4q5Kp3x4jjRdtedeWx5bqZleuVNxHtHb5YOkmC9hWRn24FSEhMjI/
CoAE4mGSaQrL74QSolqRgMBd4ellTxWszjSiAtlvX/G285JLU2s7+BZ/grCiEWL8
kyVkofaqWNIcBWDOZrfAdFar6b1HX05LaNWCtK/qTdMMaiYJqjZMWV+iX1YKh2zU
FUkbzlPY9jbSyTq9zi8Di1OfHsQyqmXf6kzAJ7yPeGuSIMNsiaJLlHlo91TIQ7Ip
klafqpwkraUjf/iHHfv8lCEldzp/BUTLmuxAP60CtdGYFkUIrgiQCEJV4aCFd+PN
pWv4t4Q4VGsxjMRu8pVUNNDTHnJWZUHEOw6TYZSL/RacLSNEycBrSr4lEBL9FocV
qD5/CjuQtBKHSxZyphqHHtDJdoUb+GKyTGqiF9Xk29Ex6KSsbMH3KGok5YePGIou
STbJEk2pU3JbGUVPgZuwAGXTpLnCKAfLSjk6ag76RHlph2Omi95c0KU3Vxlf2XvO
dRJh/jaNZsVbcHEOHlEfQtZuf0MZQlIGUmJMVWS1YyattfWrj1EpfwSu7E2mYUFG
aTtwKspXZ4c9m4u1Spqfd2OhbBDorPchnGCeuL38THgU2MCe9ikExTO2u2cCiEZM
P2RuTSDv/TQRQPsrr10MQyQgWqW5KjF/gC7huSmXmJb2IQ827rFmSmNeU+gW8Hwe
Wm/0FzNPTPh9HkFlZkwALdooO9CI3ROrjsLrncobE+y0Ly1SN4vqHmMxIM+cR9Bk
rsguNkbhShm8YEhbBEga4iOrY0ZKl+gKwEzV+SjkXBsFgXUrRbXjcGc1w+JfbdPF
+fbFWAObOtSi9akyy/cMJES7pufcCVTcIJLD13eGamFVpnS6QLRy09meCsiORs96
MDsx3YSpKPOAoh+DdXriFXu3YXZbXorAIwLz2mtMGE4KDwM7+pwEAylezd2+xLIU
+cIOI5jcaaxZij4i152x+cWwiApDWPM8p9zKXBq29KsgnjSY5PNfSxT/m1EGfNLg
v1HMQMMjp1QaQ53LyPyLXcq1MpWYHeQIqMmRS8T9N6B6hGYd5zRfeFfXrt+GYXFI
7frXtP5p84hIyy40o0KTKtQL0z6eLDK0Atw03FQpSL2m24FdQ0Vq9OSl1UDDJSUE
Rbs7WexbOFBK15enZ3CDf4GatDTDcZhRs+wO4jHqkGfN9H032MKtNZzmqcMbn5Z+
5XlkuzO68Sfstyi0WHmGIO9ZaF8FXDVWUkUAOb9JXwyickDrGRpcCIHokQLKm6j5
7aEo5e6bSAKf9FV+m3RXRKJvRfLDZMdEj0UHmlK0RQ/vMBdGr/95eU5ShvYGlZkb
fx43dZfC/utGFLgSZseVDoaB755mXmnO1ULaDO5Y1557TLI052++0/zgTNZmijuu
PVUyr4Vo9sIXMMpkRosAQclIn7s8tw1sRrW/HyPBG8TM9Yt6bz+rvaIhccXz/RSX
PRB8lUOJLAwVaB3fA3CgDbwyuSvD/n5kNyUhgrPFtcDcyENmptSvwKBa4m7twaps
Uk+6EIzbgywnSbbuvCuCvbvD9+4moe0G1+WIeey9xnk58IZsVCfn0RuhD4pQx7t/
N8TtIcWidTaVq2mXXINDE8zb3ls51hJOFnzTKGHr0LeKCS5kzPajp+hSwvFtrCOB
9I/E0gzSvbK2s4zR66ZIXLENuv/DKbpkBlmxjY2kdOiq2HUsOJ9O013e8oy1mIki
iL9/BgECQFKqYlvGQJJ4uyqs2C7HY4VJzv0YPRljD7xvyFjMcjyNnD8j4/cDMDv1
FSUW4UhNgBO94lTzlGFqR4zxm9bfTd+KjOBl5kO5cjs4ui4ZAkebJD8AJBzXSSaL
+5LvqoXUUrx9S1d7q3ONbLct593nK4hDwAqCNTaxS7J6ZT/OE05DaaW8tRRK3KRb
wworOz+2jpL0qFTXo4qu0d4KxYZ7CamCbhYq36ghSzzS0v5d5WMBRlozv2nmaIbG
T0BSx3yt/ABYPbuc7D2KJNO1ratBC5I5nrPNHlk8DnImNdR3yQKrlhpl9FLGMTi0
0R0Ry4EdOZYUXUe6mDz+Vdg009pjbQu0UJeP5isMq3FMSbMa96Dd7qSMGUsViSdT
aPzYYGrMg82tBOsyrhWitD3UUNALUqpFkTZcQBygWXAxhlEjN6QLoc11Q4HQiTmH
qdFQ834ngjola/bQlE1sknZsD82OiGbZ1JyxbTYb7Rd3yFewHffnllJtl/o3gopK
V/j3rhWE0CCJGSRZ1NXY+E7VmdW6ZJ6zWBO3ndEb0iwA3TgcwlcfoB376w4uyqnK
7a9pO2beRIGXjfnD+qWGHTxSEU7T1qapZtdTdnqaBghCELSMVW1XKqIkh25rR4HM
p0QTpChd0MMJmLI2wlUfjOE9JO2o3nu68AFkc4B0QuFTRY2hiFNfBicHBCRO7A4Z
5SqduHMSEZYjT219vGV8iMLjFsA76hbH5POUtZPPRoVKWE01fRqv1qq74uDVY/uU
AjBhTAajXopShvsvuMBgEWis3VDGHKJikCK0Zo+GavnS38Ysi/TJOZsYnQQ82foN
DKMEQgU+QMUhfKqfhfuNMwSL8nCJr5olwbeBeKWUjbEUx8k22OOou1ausSkMgLGN
NvlAMWNQMhh0Zt+OJxPjUdJ/WUiircgngxzWzlzN4fZ54vftpBdg4yOI46kWXsvr
CJ/x2+Pd5hYXossER4g2yN8XXjHUIj4XzvJpL3ByHxpfz4guJVrZVePm06TSVPLy
V6xdbsefu7UhzFjpGVvgDBBdcUs19WBQNALdsfCEZVRk4KQzGrfL3GE2JTF7zhuy
Zm7PC8OSsR5nR5VuaEvrDMC+8iDam74rY9osV+CRGEy8Y6VoV3KL396GppmvkYdl
SQ1b7yAflWZorZn9Wz9mKrIqNtEGGR5wkZ/jn2CydHSpaDZSJLRxyqXB3EbJVPlv
vNhPzrfWX9QGMbN6WjOAJkohWjkPviAEzxVKWaDDJl2jepEUpbTmhl7iFtkrCD+n
Xnx+ZVhjwq0AMukoMaMvi9/RV++HDGAH7eNkqQXXwrDKYXq/KBxxWFSFWRoh/Lu+
jsClm1987LBg2pdVZ4KgF1cuRmuFbtzosYMpjEnThxcsuPoXFuFbgnfWoFa3VG9u
i86lwmNM2g6GU4kCHChNzvD7SNXl0MW6j1VC5F1ipMP8vV6UV0kODGZFke8hzipG
QVbg0wRuFyn2Jl0QUhhmus78xxDvKOER9jU/BCZ3uxPoJKQnJ8CxwajCrFMkOpFJ
rLUsnkaD9Rw5KreD7BCBBpadtHtM9e/qjzGbIfVknI08Wcs1qqKyVqVnSTdPpyKF
vSyp9VnWyY2F9hGpgfF3/KNGwfB23hwmNNxEmUKRSIigfWSLTF4HAqXJgr+kN3Wn
dWAKWyZhHbgSxuhiZKJh7tLnCzOhHER4j1fx2e9leEY4YIq+QHVdFggU4Jo4R4b8
gCdvjkbHsAcGBYpVDbY5I1CwtUrkyM42BwDa41cvXQcHWPA5hGLzRbtYFXeqLr2l
bzHdZ9+YbKygSxZdiqyelDIf2VKIr4WJtG5lk6hSs4QXp31vV28Vxx0ckFBZlq+m
6a69VWncGdUEWSaYTGUHuIuYVdqL97PYUHTQTMYR+ldiqQeeGdSZROMxDL+6R2Ow
cdsqE1/k/QP1Cio11ERYSgITHpFjt6dMW3YGriyutJ3KkyKQ/bBYDZiYSSD2yf2M
wd9unSsVC+1CmA1ftZLTLrs1evV2eoyLmf66b3sT9RvoY1Smk+YCinnpbvWvh4Cn
4PKl7tUxUdVKPHMFl7PnN6ezqEOMN0B4jRGRCLkjKL3MYDWCtb7p6FBMRvEcaCYw
DOvi2G7x3DCqNdg7pRJ0ZKixiEyimMOW4Riw8aSt5T+lF/uhjGmp1/VqGwYmobW2
k3TXUorPp1I8N69eUxBi1k359GSxT5OvRhnSGj69ZIPick75NCCF8NPWBY1v29RG
9YNpJ6O5k+dL60eMquyTTY/arBXE4U4WDSYVSGJT0q60CPIZ2OvGOGHceofrQIP2
QPRRiQga5o9d7mZxp1EspModfRLF4lrIqe0stL6MguBChaIy45fTWH8DrLYyQLud
YH5F1AmlKLh+a3Afks8swBn8r5VRF9APU0Y392BiYlquCorjcLmOJF6ezoJIYcfv
6R9yvW5a6+XoT1btvFsgkBdxExllvcdMZjPdCBJla4La6IBurqLIZR0inoFyYw2V
S+PvemU+vO1Hf6P8mdfu26Z95j+4/zBbfURvghI9HF2XjDOpL7gT7fZhCXZQNrrZ
G/Ay2BTR3LCcNUVSmazxQ+1y3ZM9wk5APpURX3gZ4MWPI07sIkeJQ4NKpa/0As0Q
Iwc7VB8s48Kwduqh80ySzj69MBIfNTxGOdoja6aYUzxOkaleOSmSi1+OBnPwKFfD
4YfIwJM2jR5OkSXVr4Ba0sTcqQ9V4ePn4Rp1pg4a0CEM3TrlXSnVw9SCnIz4DSkA
5xY5P94RajSkBARB7uUikzHaqWnw3JC0sq/ihu17j0oB1Z6PyfTL6Id7fnst4WCD
aImvREJhLUO0Rv4LeFX6e/LdFVBHhC67lgqFxv9LmOZu21apUACPj9hdZLqtMjFK
QhwbbfEK4S/teXiY17BJBbW1zPXMhvOdT7LUJe1vCuO9MB0yYOSc5lePfvhmWnHr
T5rFkWYiAvT9QeGiHikb4ei7w7+4XEoLfOv3wDeyLEdqLKkaugx9pMQ6JMw1r9RA
uz15BHnS0tKJWv01MXigbffZrrB8PPF5X9njJvyY7C7a6E35KiwnkTfL5/v6CMTG
2JZFdm6id5yiTL90WDtpveBfBSKccBhYpeT7Pf/cNdIntlAmytMMtxNlPWAiEknu
N1aaCJbSeggulp/sA86BkwZo/lz938AqRzTk+qXL2VJxIFjb/C3AojutlA25/Crd
01i5E/dcO/DzNibsuyALg6URPm+uroh++uaI92RsLSzwfsKOiAvfIELnqvWwXpxJ
wwFIYqNlTYn6JwVkr31QCGoLj4h7seOr3+cXk3NNw+7aMC8ZwJqa2BcxqQga43KW
NqGXeAUG+FzAcA8WREemazJe8t+CHOAXtFsFv5W0r2Adz9SAdzQsUI51itcjjwTh
/P0RdUKzTL9SQguGPCzzM8U3gPXPiCuc9cP4qiwc2YkLPBM2vEyJPRuhgdCJrCH7
gYEkSXXTOjj0nnfBJwRZh59FZFCsKnEBNeF4Wj6nBfT90owCeI+lPTGxLNyw++3v
fjR512EhbDfGjV0/YzfNlVs5MSxy1sZ2TwRhMIjTShFuV7JF7cJ1ouULsiEDMgbX
6+/P41ufuhG+Vc/FlDFT0+KdW5RyBj+UdWPl4DJ84M9lh9kQjV3xKIaG3hjv03ny
ltmnrN/9YXvwYg4UWYO/R74eyEc5jukY5DfYVUe9KrguBhwiZmEmz/SHJidwHPot
vO9+/BiybfaFoQ0SaYYxUskAf4DcHkd199wgZA44iY2Ns/HKjyhJ7c4uRR2uROhI
4OSkIG2QUE8ikFlRoCqqxWy4pb4J+Qs8iLAxjxxIMEAOSRFaFJo7rU6uG3zRzTTR
eoxJaUVTVJqEJUKFtFiuPqrGOrZjbf+zRIXrjuFDrBmSfxdeoeKAKANWLTcVbi7x
ar6/EI9ySBgaqIpI1zK8Hyjmejp9FV7fwO3Ln3IS3qEqZU+XgcyauvRcsRS751yu
hp2gjsKUC6bFy7nBfOm5PXVB9ZNdpJureBrgZeVOYdUO8RL5opYTL8DXWw30FDZq
7t0x3ftHysvUuZmVeG9ubgoG+ropaGVgBtXcew8Tll8b7ukhRy2+vD25Luca4GXJ
KdfQQyqt7OjYM2rFYfXbv+cyqLehNUkwy5vCCTKwJWQZMWvz7KFGr/K82zR+EAN/
VUngnevA0xaYodION9dceDJiy5HfU7lfdczsziSRR+AqZeQXqUuEMgZEB1CTUInx
KNDgPMX4q0f0AVlebML7+JgNf9lIfoxg04AH6QlThd1W3OjpzFfWB+GO13DhTvTy
XppPlIENNrF7t1FcHeozffP3vnWY6GyBueFDEDvxks71pTXerpqoHxnEfRuH85l/
hbcPdgB8XEcNv9kyHfr2zB+ZCbkJricOTjkm40G4lZOyfCLI7N9dL6Qk5KiyJ+Aw
eX2vOQCsm1wGjOi+UerhoxSbZ7U+Cxjf7mKbd+Xd7AXFj8XOFp/ryLgMPsxueG9r
7fpO1CuPSm9r+I7iUkwjxsYf5old4t9WiLlUZ2VfGaGwFwTpvYGwLVwu183jm1/j
Mp+U5dOkyOuZ7XUmqd4yBTMglrjQd8mY1hsd3iA5UMMAAqZq68PbYU5yOi94i2zi
kbzqLdDGbsP3wU/+x9YNFN8y522TN0wa6Mw2g8cElfSzU/oL8TZSLLnYxet7gWEt
t+Gx8AcuOK03qvmi9F0hkyh1HJmH8mC9e29E9j8uCyPHG4H+TMGVrYyV5+owZF1L
WA8ryClzGU3RJhsmN7F3WKI72fosV2LjnxvQ1085pGNi5mJJfyT5z1LIC/rPEA6r
Qm3HnYQkp34LOyJ9K0jOBWaNJ7YNRQadvddlz0iaDVCdtljVws1wpasELynbkpm5
1tlqTV+c8yjwwt2QCZwO5f5WxXVMM2iaHCg2l1FHj4dMzngnvIAWCtsyCVoQLkxm
PJ4h2nZfTVLgVsUTdaEbT5bBlwv9ro4yPejnxvHozomDgwt5EU8nekMwQ7tGyo69
sEM33MbiwZ0K+3uE9wEa81e9ijkIT9Sio1s2Ul/+oaS9DvhY12Wat1PIN04JEg9X
nBSh3AOB4NlGDU2TPS0DA/QAHfxHBTasfPQkfneMsTlgslnF4oaH9fRXOTFss7LF
/tgbrJfZHN/gxrHEkEsdVG7Km9tuHQeX0rJbsL7ZNkGMw6u1VRRdkZA1dogqNp2W
qIEnLxlTvITCqxpy5stUPEs83ZaG4KolUOhtap5dBg6p8eEDDT97Gai4rBPefaUl
MVflURxscMGwKLkIsI7cMmhU/ZlghDjJtdijpnF9Xiqvb/cf3I5+lxQlZpHaEJx3
FsxDJ6GDpOYjvmsrlfk2Fc57Z93k4p38TLyqohzQPT6vQL08MMTSTsIFqda/kHsJ
TJwgkqHFqtqNRefgY/AykwfBgkpuktlMwoUfEDVo73jXXPOmSfpy8ecRO2hVZkXP
T06CeombJcAFgmm/OfDY6k18vKmShgA2H8nxgg6CZ6mLKGw3kt/T3HVFWbtzN73c
hjJQ80DDPDVpAhs0FbP4xfQ5fezQY4/bU1TClPfvZIhTGBPK+4ej52t6trT+5yiA
+7fkhp0V1J5QzGo6G2ZI+a08cbD5ipFA3FVRavcPX49BmDeS/GwqZuS4A5WgBMkM
kMadvf9QvF1rzs3t2yok9uk+lZoO+xjRFpPR0dS5DrsQTfvH8EjcEzkZGK2EXJIC
ecCuOYI7xlc3zNgDCYL8+oM26+++T3UeOoQNaoWoS+DQZO1qtbHI0ufrvIlsXdL8
jE29bj29DhRQ2L1k+lfpRxItC39p9I4VU0vAQ4yqsSXB4d1HqonA1eYawQ+iG9hV
ez0WYD5jwpr1xCIcD5jfkqDpjxr0CyUqJqs4QQ/7nI+gHOs1HbppC1i31YyQOF5r
YHTcz246GklJKoduS6oKeyzbpLJf4sGR1YIk/qD/qkckkNRqMTjcIo10S7QyrVQ9
goCTKhqIsuKRloyY9dJbK1SR1Z9KpPpvHnhOVKQLY39pa+VU3nZUsPKxRD8N/q4P
Sj6nCgKgJrQcELiJEzQyy5ps3UuFyxCuYSmzRZILYoTtIn+Ov2qHDR0ZcLRgYX6d
82ZE5jO4jLMb4Z2SZ74NDvfg/EPfRkZwm/9LiYc05gVRAsxyFc5zrgrkml71ti5S
7Mc+Y5TZL7swi2iLMoxERJj7Uslsy0LAsEtNpn/L/w1AgkdBcrWMyPIyKbXIg6eW
vZ+HeAjiRoiLg3qBdUnxeAUxakmPRD59MyhKvb9RKZZfsUGtf8MyBjTtVRXabDk6
iZeRglqapgVU+YUg4F65JAEBk22yaREcEiyF0LYroyxzqHk9bRXB926uyrfZLtWl
DerHQ8pqJrqdjo0FqVnyNy9wDEQX+DTc20C5UvCOY1l5FFVLJPpOSUiASai+zOPF
AqvKrGGBQ4wBXLQzV05jL0kdUUlLtOkKCb3taRZNfSHPjSCeYyWglRkTrvbX3nj0
+twyX+oFR38jP8O3M8Rpd2GEPPEFJFH7Bqi63HgNXjaoH6XiIQA7NcGKHAv9w8Jb
N8oRyTATU/IIepuEjOukinG3Cwx244dywW/YOrEJMfc/Au4vMS41iQW0ZzHevEvm
mM13FLsvna0Lm67X1VdXmcrmDPMHntLk/TEBcbQkgztcd7MmncjP+3Fpq4RZdl8Y
uoI6fmLIbhiHnuaZhL+S6lWZJUwGGcRS1JSMcIOi5n3HXzxYkkmq8tP8HcGVv1EV
31jHwaVp0CPwa8vySA4kMKBNz00sTk8JiaaoMsPoeiaUvizznRNvX9H28JrFAMAl
2XkPX83h7AznPwz+Lu1+IaeJc3CmNg/WaTbQmItc0naEOR4QYg7VCwN0XVr9bS5Q
5gCvE4jBszc9+p840WKBkzRnGapqdG5925R3zOGoPMGvqd+pW0Y58lWmOurP8GUK
xJt1E4NzZzEIoSLaTcyyQtbN2JKfszc8x71DaN/z5xfPggmKdZNnZZSppK+OeG9D
kA4nm/K1rxhCdJkSPMdgwNtqqa8AEgu2+g2EDMpVJ2AyxlxBcNaURhcejWAihtlc
QbmygG3CnD/3JIuyVH/jTjE/PDdYCkTFpDlJbUnbx/pjpPpQrkqd+ep6TMlXGQ3v
dfYDHBUDgR2LFqXKAhn6n4x9xWb7QQka9WyPe90xQGmHMV8ujk4x9RWBle7yvXrr
YC7A/ezZ3gUjJlCoUNLTwBZ4lVWE3UXeJbV5VPM1q57r1zdk6l0uAF362la4WCub
vPxR2gIp5Qd1RxWnxAkYYG0wA5/gHNdn3DD2v2BjkIu6FGj18Rpfq2z6isIubDag
HC0S29cFmtE1DKjEi7EQs7VXF37qF3E7sLM/flwVh22mZrmCj3LQK8+kV/uLLqH0
WHpIXqaB/TRjYe2MfsA1xCYjvgbTq07nKJQKsMGDkD11M86TeRl3MPGBwAVfRXEj
y1W2sq2Idk4JTynSqBwBQvvVpJLbjm0FhKyHhPgx7u1YNYQCr3LLfhep/3uw3duk
ZsVOHaqORHCMwWcgf6u0NXSV4nqh6/FfHNTT1l8um88UQqWdJnBa4e7ZaGygqMD0
450QLB6VYZEXwzPadO16m4iObvhaoprmKhiyP9njnxoZt5FvZceG6kOG2hWExTFb
8MDKxvGW1nWRR8miTFcWg4TVKgH+ZmmKCP56gaIaUEG8fYSTdjfuvvFtiCGuF9B1
REqSskGEVQJ04XddD79/Q0aS/qft1MRz31xjzotUYuw4VhlMk1sd6nyObbnC5fQq
fPnkI5EAenX1qJ57mTrwQ+wPRehwh8N7lhtObVF4ih1r8YUxBtTLJlefMJifhFn6
q1zeyxRW0Og2fahfmj634CczGjoqFPKNRs+EwwQi5dFWdFuyfqy1NievPtXLDdN5
Hur77u8m9esw8Zx+STou0uizsCIoO87c9JpVHloQn1JJs3jk911pqTpDxSvmfNXH
n03Xvd6Gsz4H5AZbGSXSizTUQW8ZlFmkNQkiCVp0QwKgRDPbisd7rXTWM5HDfi2X
oMQhjXkwQ8+Kyx6AMFfbNas741Dd4f2SH1WG+J9svttfG4tUwM7mVn/hGs3k1g+n
Nfi5HshMP0dXt6uTyYPEK69HFmlPKw5cjmq3inJzAn9s09KEMqO1XRyayTNNFCJK
V11zTK58Z08XdhtHt0IJHMq76umwOTcl7puT5q2Bw7ZRs+I4htFCa+4j3Qqswt4u
F8e1x6dpnlPPM/32dsKwA70yyZXMPswzkttVT+H4lRwLSC/gq4OxDnvsVP6ju1j/
OPbz6Uikum5sxCz1RTAGtL5gcuHF1IoObXvsWpAPJQ4+CdSKgl1ubrbP1HFHq1ar
+ZND6sYZ/NV4NM0JdISat9GiBhioBSHVXdutnl+lEVv0MIBVstqZIPV1bPif7Qms
OMsDtmpqNkbicBUkongfHDkFszgTFnwp0oJF3JnBxJm8+njsQlp4xI3gLwiZjG/g
aUsF93a6ZCT23Oy9OFNf3ADrG28FvgVnqw0dDCWFRbsY3K+fdD6MLA5pAhY3JcRZ
kb9F+ndgf7llBbTfToW7issjK4Vm8stbifMlOcOMc8PFDG7YDCXGxE5BpB7LoRyY
a68zL1bMtzwLmn4/wo3hTn4DbrvTSGqOfI/5VJI9j2sFoiWHOTJfmsHReTCU/OWH
EaaGyzESvoPj2t1xR5c07Z0jY/fUV8jQtICzBx8THYf8MybfFQShIYmRkbprP69v
mBZS4snumhsK8rVYTt0hNJVsQe/FSmltUyr9EVCLLHTVzlYybp0bNmNaUlkscgfw
X9QZgZyYR+niRIbQVbDsFBpLNj1V4qFMB07y0j1jQW7naLbffZ4Lw4GuLYSh3159
BQowyTUi7J/V8Vuoq4/d5UybOHvMJiFkWQIENSb1bnbXRiJ0pwohUeD1hy48s3I4
yyI98w5FnxXpzcQNVMoJ7vExX+8LK+k15u8A/Se1a80JVRlu+Z1SX/kKZmS2sPxM
3ezrz17g9fBoRdhN+cIPnMpezxOX6XrgiEw1+II7q8tO7XmrVxdI5w8n5fAnENLJ
AXril7UPjYt+dJcIeKwlRsp3qZz/6FaTwCKTv3ahwkF/WGDAwIHBldSimP0urhkI
4rze2uMXtNiGPI4KcQj3cwdaFeA7oYO+Aa2yXtskX7IzQZSoKDXtU97Buyncp3VN
kqrTqaaseLYSFIZKiKNd0GcRIUeiiwLmmrmX32Ov7013xoQqbROSSlJ6iwgw4C7U
d8B/jNAtPd1fgF8zBNrV9xiG1N/Jm6xhiZFFCyXujwr4Luw1YIHUsPVmdbn4cg0c
maqwxKVqMW7hhW2YhF2waH9sif2QmOXsKhvLNav5HAO0llMwwHu4rCsf32hFjrDb
nuQuSVamX5+biaPZAxIq5j7a+vptopjxkLQc84PFRae/zBbVSz8YX5gOSLSRFhBb
a+ccUsfrY/bn/2nQ1qdsUPG8L+fbOuVf9mGlJ7eknZQLaWG8pWzNj78PcixvdZG9
3Pq6xdKVnm9RH8hdbbihVYH13mkd6hLkjjxsH00/L0Ni/cjli73oQC9I8WABTHIa
a/9UD3vc4xr8eEN3RHMf5/yYIXEJvmvRUImtqI+UPCKIJRM8p5HvCyFvuzLXYHwA
4aJBUDmdYyvBe2J49vEY3cGftq7TvvrOEJbT4nCEWFkc5/dnmHg2djCtIzhEuiT6
Kvy19zNZBc+G/XKgnGEcZkxiLnIJhHGdbUkrW4475uO4B0M9oTiZTEq+m0dGX47F
Yk5Skse14dmT8fsdsZ3XUIMM8xNtWB5y4I/vqrPV5vVCMNaB2VMi9fZRWWxsjMfe
BmOouEb9QXgcDXVjJBcgyoewLUwAB+pjZGJFImJzDBg6ZyuusfT4PXzIrkEhHkBh
jOk2mjacv2z181CrqOID3nhNPfesHkpIIY9UJZ21VG5DnMxQOZbhWQHCiE5EjAbu
PWI9lqdnv5+JC1JnMjnuXJRS06Hzx7uTswTub4d9Wb3dMMANEHOTsJ4ofBQzk5Se
IJvCk/MYhhomKB1M8ErL0GxGhFJq7Xj08DwUAqKGPmkzpQLtD2b9jHBozVeRFVO3
On89ue51/STI5dt2E2VMLLRH7QcBWpEVmMUDFSo3cYFVOWzB9aUleIPCsx9hiPeP
rPfPYzmk2dYWrQokfFoMcxyo5wI6wjP2UJExg31Qk+M34yxboX6tYlKAWfwWlLgL
PrZ/VrLogI46QNBAW7yzSVFBwlOoj7dmy6qZ6hSvignf2cQ9pWyRdQPNFjJ/pvVx
5cstzGoCGjFA9MgS1XbNveae8mbLST0+KotFtTaMkPVeQJNCDPvaiMLZlfMZkzYo
s2CvkoKYoNoyAAkq7YIa5KDg+2auz5irBI6dwQifVC4HyKq4hlnqv/yFEYgqYkZC
qibRPg7e7139PtUus3NtT5EgwElu974+f1Xo8jQqfev3NEqGW05RWMG9Cj/OxZVs
9uLUYyZLuV7tRnYHN99xsunGIvnVdOHgIfg2QCbMRF3hu2UbzAjHChbIATOQiP/y
n4B8PoDJn6azvcG2R3+9yfDjwCGB2XzoUkJXVfGd2tL5AYFc154Kvzr0P6YM1GcK
jsn7q4Bx4Y+aZWLyZbiITzCOv3nuv1LbPJU/qQNmZDpmraGf8aeumqfFtp2j+r5n
9grHPl9oHLZzSKW0yVtXI7neHqTq9zlD5aGVuFWfkn/nibsjpyl/eVpQfXo1/qBb
71BRlJhPM64m8gkl+wsEvL6MX7zQO8DE/Q0UusV/k559awYFibnTl0MCsEcMkOlC
TBNh1qrXOrOYTeG6wUpAMd/DLFRWHtL49oup2rEPlthWs6YIApanX2JVqyb7G/mx
4jZGD571lujUp04KA1wwzxywXyaaE+Om6doMCDtO/xrZalBRNxqGmnvgk51TYwTa
zll0RI1zAczI0clu8qSTPxath2Nri6+6V3lcTHXjST8JJjHFrbdkV6i02YWSqbpj
335FhJxu+Ebopvn9eHR1gjPOyj289sNc9pLD428978Fx3i/GAMO1iUvZsce5VttQ
S76WM08mxwrymRVjR2//P9ZIAoY6iW0FHQcnrYfM7pC3y9OyFq0goZmxKU9oOSTc
s5VYacoQ7F7KFOayCD8vlmBvpy4WTWDrzeTbcRdTb3B8FobEAUjtePiUy33eaoZ/
jMsHlkXmXx3146JkyLl/Plh9GUl75cqp3hoK75QiZnEWUkit7nTT5P0Pr3Ap+Kto
eAmoYln68sDFoQItX/lRkBb4odvQ1SZ9C9/bndiJkcKBaNJd0pjgnfrPpjktQPLm
irYld/FTpNPMJaVj8PHn4m5QpTO/WKlvH4YJqSgbwaiQfYql8DnSxCzcQsWmKQOy
8BH96yn9QHTt84g5gq+DGgbrozf+mODhbhU2Eo6XDS7ZUyuBNj22BjE2C2amLvTx
VHpvtEBek9E1bEkBRERE+2ZMQlVXPwNMvKlwo/ipVWvT4Ia5WJwrfhyLWgbF91HA
pPkCBGRcObaT2SNjtcOQqomx2WEQiQOF5KT4P23RmPhQg8XsNteaIsi4phXpnmil
ftvxmJSlseJ3HA+TO7oGGboTnSsZOVaHeJp48QcrC4gH0hh4mRP+TzyIdO9a0E40
HXOCHooL1vwSB3cL3c/BKzGkkuauc0tgplGOivKS1evwrYWbJn6tJ3l/DDRT/cG3
Ti/rFSD+BjIHXqA2u9KuIcOrX8jf9IB4HwGzibtdXDXzSGuTdiHZbMtAJfMIvfq0
AAh3F21yLqtIEyEE+VQl00R8uny8QXM/4TF4shQNauwJkVyESuK5Av/DEAlLNZvT
yORgGlczBZO2Kd6ZErTusCN6KdNqwf+Wb0SZU+ClYTnI4zt+DY5gwMMVuckC3T7Z
6N02jEkr8YWZOASTMpTV3sYaz/KtPELR8aIfDWD2Tb4jrtuPWNvMWzrA6E6qKPv7
TNsh0RX79jEqK9FM2T8J3DMbLlr+f+8Tk4kn4X0V+FGHEP5eL7UaBvxi6w2pR5WG
Ur28Wk+6K1bsjCxUSVvTcsi8mWubO47lz0sjH8zmgkp8Nog7Qsrgzf5SnKzpKSgB
o+ZS7Lr+kkrwsUzEQ2hzOWV4AsP50A8I2tIUS9Yb303h82HdK4wV36f3te/mzUSo
nToWR0QVIaF+pIjMieGjrQ3bHjJV9IAFs7E0KvZrN6eSrUELcfaLXlLVKSU43hcW
PQgCI1Fbzsqopne65MdJPaVUuIo5a6oL7GZE7lN5YwaSrmGyzUsPYk4z1NNE/k8M
t9YDlKrP/xTPYZFRhBGRhOUo67Ohm8AgzzifSv3ehhq+NyYeGwS8eT7TdNiQdQNK
ykgu3K1HqaxPGFh6V0dGoLON4NGnd3j7xiD9Hx2BZpvMeMGOFhR1qfwqU0T+32ic
xIDdKhr/U0UOeQPYc5PBuCCUHCgRZtkJv7k2x674U4HewR63XTCMSktxA0c5nMEm
39/zS7eSbQGeMMGjSud1MhltIYxa7/4R3xH+rw8N1zZLqEQnulYWTLwu3w/DvIP7
JcPd+RvXIXnMSOBPuBQdy/mg+32k+b0V6hlyadI1YRYtP+ZT54DkX6+dwYCWr1CG
azInuhV4cWGmxnM4dNZ66M3hfqmwS9ZS8+lHrr8v5XgjZcXBwYCnBZHQIsE7LXcv
47OJn+Kvp5PbMNtNKtEc8JM6I9F+dQzygqUKL8dkSEZt0g0dk1XdHQEGnQoSPfgN
HD5hDFpPdYMR1tQaaOgLcERsgdjR+Xqvv8mi7LcDZBWFgkNpfI1rIjownIjrmej4
2SPvHQpNgwUTlskeLXE38qheBYFVY+PB1uJrXtcuVNFFS0UoQJ+SXwLYG9Ka5fuy
ltF8NHsEt629Ib9FaDop9uSf5YNPQxUOJ4sms7Mt2smXbcxrWRN/PgLX+ER8/lHs
yHEzyONSF1BOSgQ0ZKJJvupaLfD0kRll7+SFeCz6+H+a3jVJnW0+QTRe23wLv+YQ
rNZbbv1Qd82bAC5odcBbaVMiQJgZuaWeLX6U7/vlIOTOJHO0cDYa23VVM3fmrWq9
YMMCF4jey9fAdOYnGMtUU4PqC9bzYNBmEtS1DahK2OZyoIx6RM93l+LZ5BLUEyN4
6UPBRybHMRh2EPGiEW0LezMkWOd5MsdlwNbrcpOUbZdYe9/S31oMI2OX+zvnhdbb
wToWRjo+Ty4iuWJF7IvUdzMu5l1H/AnSE/A4ISRIiPKJUx0UVKr8D1TVy0/bK+Sb
ILUC4fganEKiy/sCaBN8G5m7UPpo5aaY0V4WrnJKQsHNthtPW/iDel3UlHKYhJum
I2hrZam2N/wuP57aAPVQeQ1guCjsYD18gRbkeCQ3MND/s7v2EZ5jlvHfKe+xyUML
0fzBb5HSR1ZM7YQIEciN0eldD5yCr+BS8hBIcLRXdyGRsfFXZV1fhrjmfso8tf7E
etHz4PN59opnl+H4QMtN9fbA/E8ZpH+C2Riciqq636NTm0LApsA6B8QGgK4y4VGe
PdA1S3JyOpdWDgmhp53EkbL+DgzMJxUq7G4H79sgYHPwXld6K3+LMchOUQ0jeItS
4higNlpmw3pCCIW6yxrj4xY1r0SvHCQthbLSRk3zIBhDAaHCwaSxlZA4Y914EgEK
3WTwLJv2UCmdsrfPHhjQq9Bec4CzPi8OdK6PRm25MPo2oT8TYcE3GYPmUWhHrg33
m35dj810wQVaYqk/v7KSrnmuYXHTlnavW0FGCu8NRMtvEWRfJ/BnIq2EcnB7RJXD
k0cgy0agJvs7PwS2wz+HqTIKYDWSKDuH7XC9bkAhv9moBu+MqutvPbbVpImWbrxD
NzP6qdMAM+qC8+feTtXBM1HEGA4CHMksiMMVUX5+hFWBGTsV7Qzsh5IO6gAGokSw
LEv6T+UVdniFZwaws7iwOOYE8D1XD63CqT14EnyG2GbU1XXDvNYyuteUAAR1v9zi
4QMQ1+R38wPEUIQvF7xDrgXPnjXKy0HQI26a9m29dwhGbZuRufP/5NWhT4PW27X4
Z3PLVkI+Fg2ighqBE4X7KLMI5tk6vYO33DGDSxkJJkEUWfNDl6AAdMGLV+PqQvsW
eE6489x+xwqZypGIYblMW+m3DwgrtpoJniKAIu0ODcQmdmPSL56rj6s3JJmiDRN7
aXmWwkn/qbaSP/isNqZwhMo3+KCyTbPveoYp4R2HWZn4U5xOy/dNWcReIUda9pIv
CVfRoif439qKJ3WMkLWOLImVwMCO4vAdhsvJYHcD/iYDICPAB7WsXPO3LvEnpO3P
x94fnScbriH9tNO4+TwU6V3Z9wGE2elJ1zf4hGfeP3XcQfsqnTiXMe/9dfpM5nno
G/Ll9jEcN4OO8//2m0S98f3SL45nJ5CfrBJx7w6cHzi71ZI9/AMp885oCgGVr0yC
Cx8KE2Uy+46MYdV4QFyfwbxkZ8W099KasSVhhJe5if5UXPUFnCoCLZadpwa9I3PD
NbOX2sU153hRpDbEKQCXhUU7sqoAAIXMZpEk/kPGL4fNqckD+NVYoPPXNY446gxu
f177ssRyvuApp+T8/rMJLcTstJXYKQqNJCtQeiy5ponAQkyataY+CN7z2H5ebouJ
5+/WxhBUC26jsv8aZTJO7BsBgIuriOVCMgSaMELgFtoxYVxKkUhuQBZtWtsVVOiM
ejHAqFDDgH1hqlOHESULExTe4M5Y8/13JhpWiZWdE9M4GDEUp/WOu6MV1XPR7q9C
fnaXrMo64T0x4tLI4FyhiQ/n2PVStfoOIcJSB7yYNgyhNCKeE1H1XX+D7/OSfFGF
9g9mEi6Ch3NKqpOEPuyB/vRt59eBuVY9NldcPYZ4urHja1u7BKh45Sg7rnJ63wfU
EdiNG2fzMj+vPvOmRqVdtNAGaOGKOCucGxiu16hHanqxBolCF5vAlwmm/s0XFdR/
viJCtq9lXTKHub8Ppmu7j1a35t3DOMjJdI1BCvcJrzWcmeApYiqa3PxsNkfy7+jE
RiLa9TmczpMiQSRRAeuuM7r/LSlEodY4DpvUkLg0HZ5AcTEE/76dBvK4e3O6iYUY
Awr8f1eIYKri8DnefwUwOUrVnxVxvxC7Yf3NAB87KflQ1qX4gNqL4xwdV3lSt8Rl
VyD2xVNCgf0wCq6Ne2NRBzwd8ehxe8bIee5FhGL70GGcO2EJrsxwKL7D0eVNDCYU
rX39k/tOzchR5SYJbI9Fk35FPtOASm+FHdJzhqIFeJgE00d/QDDPrrJrknsrPLA/
klo47fA1PAXalSaKgWsO8nmmQOID+mXt6937p7nKwCe4JdVKyshBeFBqTbCPZpTz
F6RlAfCAPQaJ+2W0fCebL/dQzk+19OEhg4wTEbCJ0MsrvyKgbU/fxzZEpJNZqihm
7qrgib/RRMzWX0qFrbwjLVQGAgeumRPrJCNgBfMjwGvreaEcKbZGnRaUcHJbGb9p
rxMHgHtoT2iT08l63KSicxO6uI+aogbiPbWE/9+2ghAD5I0Y1uraqLeEw6fzyEuP
a2vSxicezDgJpOtQ3wz2UVTb+QmkTcnzKdjvDGyPo1Qt4ubLozou1vtXmAmyfC7g
ttinSg5+TLehWxBQCj2oQEZIrKkHNZMl+0+Jt8ChHbrpNSN9vc7zvghQMbCjT5RN
7WttSJORqdaEc9WN+HXfrFAAusP0NprdeJd7wnUpZRofCRYcWsox8qy1iyblRNB/
s9nt8OvgSNowQdSW4QfVbGLhx/glqYH6cKtHbzATCNZV1tY8QmVZdtlP0WKCqfjR
6cbDnzJu+hnPYIxhR3TeemG+XyaDg/Nuq09jAOdRvPcf8HnfLXiY2xvGDhHBdp9c
FeRZn+Gd0yrQRYh9PwyvBDDcPYMz2eSYleLnnbzSV5/dTvBkjG1PA6Kfq0Kmv1Vw
pkDoSnfBWWl9tMkO5D3LeZnJwXe2R9HxdKKg2AVC3L9qeHf7hzPcHC/uHNaTdbuN
XW//NsH9SEznwYnMCmUNDMUq+mBhyDundituSqpSJyQMdYgW3bzBXgbpQwXf6gaC
Uo1o4xqT2feUfARymWgBcuPtHUBdUymQPe2+S4CCKGf5/aqx8tfTVnNTsv+7y6Gw
MnMQ/TFzgXEa2VkgDBOSpX1k+DFeyU4oB0j1wk6+exZF5hwgZ0h3egQrnJUb3xKJ
Xp0EgGIO4KQdNDwryNT1b+6b85IbvYd8GEsItpWU2BCwD/M6bP3tNQRr0a/sw65/
DtYManCVMV/f+qKMav6+BlrAH2pWgGGZPEG/fxHl4rfPjUvUoCZpFjXYIPhwd6u6
eN1KnUmrUtUPAuxFVQY5QaLjBYAfavnIKzaaboN1VvVuaXL5HATSakJDmtPM6PFZ
ohL85fLG8Cc3llTcT6b2Amg8RuxLWagoJu5wv/+F+6Gd1+q5M89CPC31BwebbKjj
QFAGKja0wWpwKRUp64sG8KGRM4Rhh9LyCO5nZRdXiccANeoRmC6zZulJOppbxNeI
nBh/qv/EMK+8jYmwGvJDcobgHSzMDt02OK/p5ebeT4cjlujIcXJut3fOeGj//LTb
PkPg/BMxNQJnoVE04Z17GDKRDoGgUCxR3aQ6fAFuRTkmcKtuRIShyfeFeSOLUEZ6
GN7VShAz5YCrEn1X0ja425uWvvpopgB699zC54dCrsqErMKttsHlyyIhxowIyQ77
ELGCSLeG6EUZAWGeD5sqEjoRT+cNgAa7nlrdIX+9M82ZMG3V4N/ip8vfAB3TCKKh
l41GuXnlaSxtYVzB8eDmMr46KDnAXyXsvxALMgfaOn1/TLKpXxXDGArb7KSzgE26
6+DfYtv0M3a/WaFL64HJ7ErlmSWCSz319YZ0yFD/oDAFcb4GG2MlyYxR5ZuSpnx8
TYXC3IpCCoIs7RMpc9MbEZBhs3a98H5fATIb2Iis9oTqDFXT7DcwUPWfW54Z8Law
TUTgIeUBbKx4cPzQxG0GqGotFMGC3mvdqdW+kKDJUroyjxypXrndPGgjlCgEn9Gk
+ZrrP7V2gETrFra+D7eynDn0iG8mjLP8yiDf3prGbQrIzx6+H8iOUr+8IQ7CTATy
xoOrNaxZytkfYSrnspHvXuTqZiA16bk8kzPlb+V+z4vKe1N0p3YMSJGja+cjTTxQ
CTIKs2PqQsvtRwyPk9xi3i85SBlx4v/OgyPHgHnfWe7TsfAxKnfognpQkk615hm5
tDUIdqLGuU1tc9aaCgkAgsWZvgN8667Kty5Ldc3WW7j5p1czulzb6rSz1zX4FjmN
kg8bNMwsx0B4uEULQdC9SgRtv1Q75cv1rzcMJlGYgZZExhz0L6Juh5bvVBFTWiUZ
iL18Dfn4PEkqHiv+0sDT+a3CKmOV2u9KDau8vmXDc+/eoKTMYnA/e2mNiwwPsKmn
ynk3iqZx5RFcR6aJsAhJLbF9Ggzc9LwUk2kvhYqI/OUuUh54wouF7A12xe/iuvM3
LSiJF6o6IlTBF4PPvnQgaUygl2ZTsTm6G6K52H6/HPiJTlb1+zccP6aUWAru4Zps
b4ULqBLYeZ27i1cRHyj7RNk6ehxPy8JFDG781sG+Mj8JPc9oT5xfJswZTNuXxd+d
OfU85vjaWbKw4En72kp/thGxWMG9uWlB7tN777ABW4zKt+6Eofq9jG23Kdwfn/fA
xfhPVqb7x4Sigdkq4RzzgWthsK35gpLvmMbEy5C4mFnpoDhGyJ1xSAIO6DtVtXUw
hZH/nZxyT2Q8GJx5j7DR7QDjr3kxAzEE2xRfiGQdQgF+h2Ahy8Yxi2ZTRlslRIBJ
v8xhNfEi4lnUVVZ2xNWV72Lr6ZQ2Jvh8ocfCPE4ukvsP9FEw3UgbJ1/q7tVht+WR
ei9r3NQW4KqKi4zBZL+QIODsmWJD+vz/b559x4c7WJC9fhhSx47pQD32cWpSk9So
9RzF2oxULCH28Te5Gh+s2rDTSkZhV3cLJkGHGplgU1P29+JWtC1MlPHFzOlJz3pE
IXOpAxR64hdgkh4LDycKf1sOJ/u3h/0dPRXU48Fo7rNq4g2D9QrpDGvl66rkQReJ
hjGLVnYLlk+o3+E8aMqTnpiPm1joTvHHpAdIhXUwwigRNkgatS7zMP1ZDGyuHUCk
vJsSpg9bHXfszKcIsrqt6EBVbk5YNik04mifgHPbnQ9YgmMBb5PkS7VOfjFFsBTD
Uberwlbl7rReklNAEV7jdYqVJPldqxkQ+eS+XdOjX1lolAoNV6UuVxFRV69sMdex
dRGUGgS5G1gGl26UYUJES0wHXZuDTPA206/m+dW8K86AC8px7H5Ag/NXRVFPgCZN
9Zz9JA7cq2cPufoEdSeAJiKsghA77T9cVn+vg6rYZlT7/3xdtKARNrsHWSwJ3e2p
T/01D+fXcjVYfGnHjDJvw3h5C0+bHyVmgIRmuWhJOIYCpxjipIiVF8S+JQj4enoT
IHmyayVqika3HU89T68L6/4niMq9cm/uSUVFqgh13Zxf9dDWMU5JdqspFGZqiju+
4KHhBQezRm4tijELJF8KanF+91AnoNVx1ge0AGRGmrG9nN1j7Tn92/Pa6yMON03/
QWUFzfjeZMr7mEjUGcROfDi6/mrVOEWbvBw8/QdlzPbY6dtk9Iu0J2zAtArN5UWu
++VXuMp4j15VDKhi4jlp1yn8wQ03g1SMzC9J4fhwp9Y86gDd+WQs9oIM3BOfJmH6
jq95RCuWJe+FV8iwjMBjtKSaWrdIcEIpWDn79EhsEZPGgU2qi11AXN40OiuAeAK3
tgee4P8DToZzGT7ugYRhxapxReT4JoNSXg9zX2v6GBB/Fsch/JHPmLkH7sRTwKMw
CzyBg95H72cWaNFNCbTXRCdtdWUPGcwA2+JrJinbgJKTyrARlXv9AnxvZnOf1+jk
5JRE1yMQz1yg4tfbwl4UZmWrwKYbGfsNixmxLiBx4jQ7Qv28gzjYXAg/j9SGGArJ
fGtNS4BoYs+9EAzXVnKLFm+D4MpXblst9LDKoeywrK8l6FOijun0MZ/h3U0EMg5m
gUKKCqJo2EISzGHh3FLajjKt8qSM3l2i537XUOSY1MzlpXxF0ntmF60CVqENpVRp
Pn/1jOUl7WkToeldvnZWez90JFysreVXGbMdEOZU4kY3uCpP5MiSfu4MU/vbC+52
Yt9E7U6L6NRMoJlDx+jUeBlt7DDjd6F7SQ4WKfwXcKViYNvCSFgvKSRrtnW0JuyF
X2jh+ai6uMi8bqPVvQOKsuLZ/7Vy1+FOoOY392YtimC7wWmi163UYNS2qIraGUGP
oMSLRvAc/3U7IFKUuyxMdqpb8EZPSieTNAvvqIgOZA6TkFLyQ0vV53gNvLKjuVr6
buMbm6XTvhQEeqiKKslCXVNfkMa0j8w0tgK/Lo2HrrL9oDYg4xcxJSHOsKlqFev0
u2DINkjko+Yy3B3CpNCmccfLaupx7nCq4zP3ul5BASaB7UkesGIt2dABfmfrrSra
SdYjmNuMYlBqU26za9CAsFMfOfyiLiSvzW6OYW6kNcUuGuzlvu4lddH3dFC1rcR9
uxT1+BVwIK0segAMfT0b3L617rFeBZ9YoiBqBDzHiQXcwyW+vTGjh0UmeiEijcZj
fnZFz6xjRWqo9+qXQHNgIOuLUgqFQEr9JEd/N0bjQdb8OGJEo67nhaV+MSqPX3Jo
bmLKDHQf/9YcEpyoWfvyulVMYvKDnB0pXV+cTYksqu4DPnPK6KZUqbToLpeyH2XW
OXX/jHGOjAK2uoBckZeOmSsiSj+ARUlz4cupjWdf1Uzz2tLOuO2RjR/MIjZBr+ot
R70ZcPapYwq+cyIqE9vlgpYyYbAvAiFgvDlDys5UINfMcQ73KkiNDcfpdVCqbKdj
PspbDre3S3/byU8opgYqSDzTbHcpoXwqDWpKhwZl7Sij7PpXW5HcYuhjpm+J5I8c
M50Q3JbnJVOxFnNRUXQf+CB92QJD0h7h2wUCVCZNIijM9svQDapQ9O9U7LPMUUk0
2iwLdM4AbR8AJk4mV3j+p2SVLpjO5Uqh/Y40PtB9lHxeJD7KIqgOqHh1h+vztku6
IVjPWifDNR5Nn3DvQL9b+GLtoMZgiLLM4tKIOQ4CsptW2N7nirYBY0yrvbQq/3kH
U9FfndIgWWxqWRZfoXRJJ9xanVNJLTAhoQrRJV3yB5xXxw3PVw5m8Elp75y5qJiq
O3zwrOejeJwvZVnepc/62p5zWoqh09M8Ex5qFaynbA/Urn/17ZVftmikQPKvx+CW
vvg/S88Y6ioudZ8S+fyJBIdAE86IHgH1dOqHHH9lzXcv95/gqJWe6aHZitdoqdA7
TPX4IvzWoIit2poJM9ylEiSSu+bPwKy3Kyz4ue+xarYHAbBtCqk6eKLIxqD28+ZG
5g/+Bv5AWvnTGJ5ahFwQPmkwCfZhbVPbr2mL1HVBkrHQ7f8vu4pNU+LTQdJnKk1T
DCSrPFdUr15eKrwjFyb5QYIGy3dQR+QvLPK/V1VGjKz8SPKGLpd5jVHJthRb+nyU
WzrB5KeoUqIV0TKp4Su8PcXBbC72jjZ6Nt7+Zmq5CcLxda7I5Ryp/rN5yNBb8AdA
RkP8VLhvbDhAH++XegPMewD34O/W9t97dIRoy1lUxVebi0XzdCMI8Ih0cSJTnK8T
zHbumswapeEnOd0YHVfWe/P8f5RPl6BHUGCM3ztpzRbqxdZofK3vsVcS9pRC7Yeg
U2zu4OapD61+VaBXdGgGFGy3fntQ7VJfOprWFVC9h3kgctNS9IhyDR5xv5tHSODm
8n1Mmf+bI/pDFGQRBxqG7VZBOraJTV+b8GcIttTKkYuh+/ZlL+2bw8m8zJbeg/Cp
1F52q20By+kQwy3pnOWWzph2TdMHArNDFKMGiv4kQaWiemDArLkAHCb7cpDBOjB2
HDYvr/MZclcCIrCOywW68JTQ9yXDBw5lgm0gj2OvE9FiAwMUxMpxqJFtlcrfbOQF
kPpDavYIRWGc7B/1LLoFH/FyS1uhs0rsFj0vDXS5HPTpA37stPQKZFcB1LqnUqDq
J/AnD/KR7THaU/DKw8sDl7VGF7XzM/Ce8NbBya3kUKd5QeBawu7wic3/0D0Z1baW
IJxsYziSd1pckN1oX7ppoeRKTRTsryLBC61vYT4bQX/SFCjGeU9Go6dcTxecd/P4
SvwUZV2DFfWyAwNFQ+XZIs8xDP/HpEp5oeU0e2Ypq2XjaIN2QpWeFy/4otqhg6ea
hbVyD+eg1dMUTFG2Gfd60ZDu2irxNAqQeJdtgSNr0w+7BvZ0tjdzpGHiqdZAzqcS
5pOUo8U7hwN/GFZZyAT9Yh635dHSXSSZCSReCNj7w3qqdHce3PPggntEQvhriwMM
MtM5fQaH9J3K+jQqX2fcEUefn50kYZebekjqBcM+HIpPRHsCjcOJAzyb39N/4wrn
NbfBu1xUGxq8yo/D3We5hWg05LX0Z9QDCOQNUMq43luAc2CKeWzoOtsYQ8RLt2zX
CLjqJfQiwcDq2cUUf8OdZ7PvQ1Mrfjs8BIPrt8GMoOardWu6LF1qDVTst4t7efsE
WGM0rilqVsFEJUFa3SzbIClRnmQiPGk207R6OQzJ546LDNvYmHD8quW71g92ZR2R
By2A1tpRkbYYfGTT8AZ/tVOXhfFTAB7BCWpRGudQ4VwomxYcV6HYDQd70LEFzIxq
og+Qi35L3p5dr3PIgpGpSmIzxyER3V06JlgnyY0UifpTsSx8jbzvtNKZIA7EkK+K
bzyCqW4ixxM2ddLZPyLLG1jFTUa1OVff5xw4y1OAvW9GDrwo45L6Q9Boohpm35yF
9Eu20eYOb4H20nheXbGg+Ahbd7gi5MEgPTzjp4cDouMD7C4AQxpuT3hUkPzzl5G8
QgCuRoaS+Y0bDdITlJdYLeBQ6DvbCsSK2JJ9Kmg9X5lMH3JYn9si8KftaMxSu1GL
U9za8wkMMZhEx8/qHySx0Tp8N5fgERidCzyofhx8lxIZkPTv66LaYpMRfgvJfA1b
qOKB8Rx3kIjPqt6DmPIqnNckjGaChD/Rl/l7ZXRmQwcj4wchlFvSHlcauFnSLSdN
3Dh1zzpqBAjbqxn5oL6TYqG7FaMCgzz1JoN1ru6bJLRMEPrEU/ppPzABkrI9ywFD
53Drr6vc/Q8kYh91IUa1vsBBtbN7XcGfg9/w7PiqdBokMCeFMl4BohtZHG5AdJx8
feTJX8K+fIw4TT4+7jdgMy2Pim4TdptlpZ+vo9BSkqmcy9uAKJPyM5OeOJWetIvH
69x7bUvP+/A1qxu2dP5N5twgGflRkDX+F+y9BzK4sN7hnPMs7AMWOE4HGEszImvl
xnsvJQZXcm9GQ819kvX7xBOnZ4UiclmYAytFdEeqtx4dqBFJ9oNMiIOrMpNmrsRQ
ZslxeEfPwDthc2R4mgWXYLgHE7uUOLwKCihF5wQkIo2NoB8AJ/sEWB8Jvt1WjGSA
3Cr+9Zc9zaGunSYE4FqHZUBm8L6dKQmGZvbTnKwDtAPdCMhUepPy2oW8MJDKRdyK
Jrc8RB35vQxMT/RjYxrtKPQ4czeAnHjw+Ov1MnDhgjZ9oQfkWDyEKeiqxx9gfDS/
9qPJp6r1FudtRe25VmX+8bipuRUYH44v4Q1phznSZy9h5nsD3nEzWGdeqhWRBcfM
YJqUo5hxDr5hu9h3PGVdD2DPUefgQFzhk8ZQTpyvc7/JhvzPqni2vC18lZI2FOdb
kkItWvQteADyGqgGI29S72K1Uo1Z+M+GsQQcO8neWMIoDcW4DVyMRCZsyI0TxH5N
VSahHpy79gm9VcoK+YGJPI2rYpmVvfSCsdbg7y8hQ0jr3cXocNHgR2hZJ1YUQ9NJ
YuoMTGcaix+tjYG54qS2+jgcw8puduclpalyu43Pvb+B0QD6lrsMKkerl6T3r5An
2rAAobyzPNwEO5Jxm+WFEX0u0v04oAZqAmu0SRq6h9fP8EqC73TMTS3lIzt76vn0
X+Fc7Svw6+SR++j29JrYCJC+ysgmy/OalRR6rb7QMgCz+ZW5nNIQpzUgiM8CHz1A
LKx5G9jm+Q5kzFRhASAymJCzbGe6M/geWtUVtPCROjeax0Se6YocOiRcWggmT0XR
paxW4Vw3fUp61etgqSR+MxP0vQnnDSJrb2XcT8ErsWDl/iXPyxJCYhmGsDiwa8w9
j0OLJ5y0mwiafabK4xycA+kxxxDSBET3OaMZoJk8OeX8WTwqmym0a3oPqI1zVhSf
/UQif2zNejV2PsW0LcWhyYIsnXECkDTgegynzShXf5zj3hWjS0qz6OsEvqTfzfY1
4x5hyz6JRZ8Ag+nt01Tvp2TqOoGVxxeATPb1QOghQdW7jYKSOLZVxOWSfTxuIfYX
IgqA+PMHV5DqVljFdW72qwCYCnsyWRflYco5dMeBW9UmjpX6AbQZ/Mgnv58wi0Ju
f0OZhgpUS+zvqwEI5lAgaE3tdxz1ty2sCOTMz56zPPyhVySxdS3XybUZE9E6lAA6
Lp4t8yUr8/RgzP8yuN7iv7280pJAo7kNf+l+h793RuUvkPsUkxid4HW/82s9upLA
w/PrsK/xWrzZlAhTI4dK2Kjb83VlfeVRN5Fxf4CaZ2GztVy6OPxCuhwk434Zjgr6
jZVLkSKKMNcDIo0tRWuYg0+ChOMcDifk0ZQERzDbTW/swBGrxDF1n/AxINbPlXGG
xglyhFVyD3DXfdi+uysELQoNbrs5VvxHfqvKlzeCoBu1U8MC1JB6u/auiHcEz0By
NJyP6wiNvs/9L3Jl+hbO8SzgvKrcLmuZ8JnOk3EMBzACU5S10jCWCt2dIvQYdyMf
PyzTw+8wPtu0waDi25AOFtPpDG47KEccSAv1Zl/NxHaChlpeLv23Ch2+zehWLJn5
ZYLJlB1XJKA2E2hOZ3iVc46qg2+mGWUteIaT5SiAd5dnzLwluWFEftFPxQYOjiJc
KvE98PzWnc+kSmwBeTrVphCQxKWl2bO1N1AGOazJlydfIOOeWZYLZ6vnP3Ig+1zh
OJbQO1mogIU/eX/4ugIbCPluqG1b16ksbG5cxL8Mnoc+k06QA/jCgxkFHyfBf2Kz
8O+ifcQRVAwxScH3wzqUnjxTfEYn0cF5b5w3tnRyVP01zxD0ReHacwM+QYFXZm/Q
HIjS3UgWaye/OU2r1d0FAHbKCFVcSx6KdgMg09/Oc18+kMcFI09bGsgg1PqS1/ZZ
pXgDfGruVSsI3pkEFsC9adz26rdL/3LzgNiKAPP3Hn1WAAfFeKOM/RADTxGqYqc5
5bUpnfr9XkPCLsGyiFZGE/ZuJQghBxzsR/BOFXae4toTU/+F+S46eVUGiuqvTHp5
CilMRmYVg4T8LIaanTVmc1HESsY6fVKkttLZEyNpZl+p69EYMudK1h4CM+o2yx8W
LJyBPSpZOvlfbHxS5SCW7+f5C81scTNGT8R+x49XHufy9vi8T81hxzFeeeo3dDgQ
0ZZPrgjWyF9hG5NV0uVitxGZWxB+zkfsSWpPLxWC+OYhUq1rk/vXmG20XAl6tEjF
X9hN7VdSPM6teOS3b1Kxs3sp3vKmeTcy8WJGi430WuzEoTPTUGD0BoEVF6U9U9hb
n/5G2uZ49zmjY8BghvxF+U2xO+v1GqfqyaL5NRCxn3FhtWGwXJy4yHN1APZMVo9e
NtDy2IhtmrFYSKmCjcwX6PXTjZplcnXWwdRUpXosslF9N7Uxi/3OMM4BSEWFz45C
s2H9LNWu2G4rf/Lonveto2ihvXTFyxKKK+4yhzt2frbqRb0rXX4pRjpWOzJPfBP9
1i1rSlj8ibc6l6y40C8/ECFmO41981oqhkFoq7HXsxSSMiTDYAVmG4N3h2hkrqCY
YpNpmHLkXhf341xeKRhZQJF9tIsmJyDwm9msiRnUsoI/PHty0qHO/njuw2rFr+zn
WBoyPXWAnrgc0WPML/M9fXzYSmaGIRg2b3J2vE/holqal591yMpDtu89m+Xxw/zL
JBenSLyr42nj/y202JeE1JRdxjG5Uqq09/am3wwHCJD+DPEOQhX3BcjqEcd9Waqw
abO1R+SaXxgAvf2Q9l5kkCmeG02lB40p7w4ak1rKglX6t/Bc06g96EdvxZ3oTYbh
2f4CDcL44U35myZE8OLlaJew+nKiDxER8UhKOl6X0qlamMYCISZcAaqz5Zq4AQbo
BZg08IiAfZSivDzCfp69DHoHQPe6vi/wvAtXPUEuwn97A0FQjYtTmAnk0EupSH4t
bH05+zcVs0hVhZNOawXzodsQam5ZLbh4RZhPMk9r7mwaiXnzS7541AEtrM12P0xf
NM9m3Bk8/as6PBwJf6N1w3T/vC/z94FzwXOjkcGaZvL9zWMypr1kypwyB+CDBpH+
awkWo+IuJPNMw+5pGkqdBzCgwQUDjSynzK22jvxzrjbUS65o3cgzezb5JBHcfdk/
+jpDbNSmybd9Iwz6pM1Z1+b6hsukXx40uoGua+G/dpKrvgKGMoL572yxITJchL/U
OOyJic8NLShzEwEjeufXVTAep/YJkSkGnUSjKqq1Py42+470H74PWmQM6vzIUfVi
CxdbXPR27F4JYpyYLvTsjSRVaDX/cbJpMxI/wvY3JU0jxEYXmmIdPCjKMoKbDGLS
kP79wETh03IXFkglfR7dTlgReqtONPh+kytY9MK8HVzK0NSjJIY564HnPdSzdkot
6XREvInpsobeHCjVFdeTKKeMCdnhJl4sZSNoPg9I/AcWzzt5jB5FMF0J0+Chw4OQ
A5737d+eIpy+ot6YGQFW6F+8I+htSk9n0tGWa/T6w7XMVP718crJzu2tFRIifwj6
wgIZx7G56pWWHf+DoyNEuTLOIRLHgZr6EaeToEBQjwHIEBOitrx0l+mol8BCVHXu
YgMBXEC73GAbC3lDf6VUtGBzoErxuIQR1Nfn56hI8ca2a2jd2honrDw6h6TMPTEQ
pC5uNf+8CvXat2SvZ+o5LBTd1GQqKYhYHy3wlW3mMOT10kMPKeI4f5F4FRnXbWoV
Txf5WUekRkTpOy6az9DUPeflZJiBt2RQz0IIpM/XFGIQ6SugcbvtWMOyqMb29gE9
FGiZ9fRXL8dabDfQ/xiGvjohWPoAkryDShPyFkdhvS9O9Dd8d2e743wuVsd1eYDk
7FeJBOK2Bzt4MjOrOb4W7S1zrZ0bRJOlKk7aPWo62PVAqDJ9Oh9Zo8hZ8YPby+r7
Ci2QayJnt2QQLa/Rd8VryZ3r4/mR06GbKDcYYpzDFAkhXWId0McdmwuAY3skD0nn
mPUsvBjZyD/QN/Lqso2Liw/MD6Lq7F2f0kgq6Lu+KpwKR5xYn95+1u+3+c2TDQ8I
ZrA4ALg08YhY3O9zDNklohXJmlGVy1SA7zUvPGEZXcC+y4imLlB+pfc8HsJ9hzxz
L6CSUt6UAgq4zCWSgWdh8Y66CE6MnJetp5XxBENcVWLUUAyB0r0OkIcMpBWUNL5l
KTlaARMcawOrHo9YUbZTuGjTe24F6DlGeqi7uFcs3Vo1jLCUx4w+q9lmxKSYsvNC
RBMqnur2DGHwGmCPCs4tqG482jK4r68tkfFYyUJ/lNrtoRI8bXlrJ/LmBprxjCzo
Ixo9nhugSKw8pUo4FbHbSgv2WfxiaAHCoXUz4lzH/4prPu474FBxmPmfIl5jpaf8
vKf9Jqpc3hcf23HU4qWoL/TSXnTIA3eSVcteFJkoSzyr9Ij/Q3sjfVXDsRy6TCoO
sluvIPMc/DOyny6TOOrBUQ3yo4C8qT0S4EWxKkj2v3+REsZ0/EpV/TRrYQkzpELa
sj9UTCwIHP0Tm8dazJW7IzFL7Y7VvzEXpPmqyEcVxhkpT0KggLUQvoN3wMVrZ6VT
HWFyVZ/hh9OvtI/ey4EOiFUknhWzmpBJaMcWNXjdSGBdsi0cJXPYpE5R7jiHweTe
gI8+qpHth9Js8kLmO0aQGFTq8wH2ad6dg2i9+ZMj/COPM45i/aFZ4li/Pcl2MErV
S3Ggtl8QfudzLes5Vgri6rYbODI6m2VxPVcgM19ipZep32aFWShjQtLBN9NMDzeF
rUgERn5Joc6Xlp5Od3rj6CZY2vJRKGLjl/Sl5Uh1sHOxDWYXRXY6hR/pO9TH/lUZ
38koLk2ahC549KDaNvfQxgPWGmlIuGWjMnTn94q4vTsVvSctJlnpVbJ40wTs/VuA
h3mFP3rRtdVrU8AqxrkJhW6uZ9lANojGWJOYabnRHly5QYenrShCwQVhRw/B0gHh
tFTGQ9dac2vvWm+VTCgoXPVYLVlmpThJAyC73EjXJGijOqnxkDcYSmj7E8QQG4jA
B8tyMbxloOWcNFnnkaICCSs7sqAvzSO/d+nl4JnvtR1LDAK87kErpn6tyblH0Pco
5mX+YzQhcTY/NhF/FwwG36WKju4TP09HtU3bvQf+w6Q+a68jSOeGPhSo2+IXRyX6
8FWoOtoTOI9drRN2iLnYl2hSn3jZi1U0daLd7XEfI6KY6iOSlABZmccF5MBwcDnQ
UQCYb/ZPILeIGfg38BXVy4Uh0F1X3N7OyUbNZ2dYx5mvQgZQsBsYCZIAjjluq48q
Y0T4xRm6vED26iiE/tskHkswocqG3OLdyKIF0jKxWsKx25nIhBkYnTCZJrIHzTs2
83731ORdinkRL1l+Q++AE9pzeXG+0pKiL7SVZUFRz3tSGq7dFkzOLHgzVz8YOG1L
nww7esRfHYO/uTd6Fgv4hsje6G9AxwRPKIjwP+A/4GD9VEUVpXi2vjjs1zUQXX1U
ZsX9055yG9fPBViS4zXmOAtnRA38H8KTEBYSbiPYqW+m9dQtbK6PKhZTMgU20Rs6
Ik2sepNytogrRTIY6YZO1XVUmrSVo7uIdvtWLHgv0jR3zPiIkUe8xMM1bhs/JFi5
1hFfF2hHfOADMU7C5jYOGD5Q6CX6rOv3JytMHAbkb38wiPOe7fNGYaXtZeiwwSiX
XBFFBdI/XTmJwJTOpY6yhU138ChduKWZLCR7vvf19czd/EaIXpAKX2NH6DGXQ6n/
sWC41P2za7Zw5POakg0anhjginT+sk4IZgju9Ka0n3q/k4JPh7QMMjQaKxeoEDrX
00jmYxrzKMZoZTmW3L+w1+HC7ktGDgE9sazeE7QAteKGsno7wwaqtOrBwOXhHN8G
UJhr3/+O6YLnDwG0rNy9Xm1QTHUu8GfbjMoizBlruGMk0ymzDgITH/ISyw7BZzdL
ZIFy6xVUqN3ajSyCPkEebJDNWmlvIO69C1+Bk7zzkHOlCDPhoqntDI+Njzpv0MUU
9FbHjVmLHt05UVA/XdgeOy3/szwVCdPBUCM6CFt+iwxNjrSeXDEcCIDLNi/qRz1T
jXxcsvRqY1XloltT9cVWwZlEc9B0Ngv4UqLXt3bC24Psy949CbWQkUcNX8Jo2cyn
LxKkzib4H9Cd8vilOrPR6LjsjECdBYEDmqUprM9+0+oe34sXv9GpCnQHlRDf+Ulm
Pi1VQ1aIUppYgihmYWV3ed0+JLwL6hyaNDIWr4x35FEdMtbCc+cXxHD57rVoX980
iHOHJ7FCSSEjWzX5LfFtrcWjS5puHrLgfZdGizi5VP6CvV7cfU34NG/5py+CZGm9
ubA6akXCkRnojflH8Z5RetolYHJV9HLs912B2P5oRJDCpkEjKLnNZZfmJ5csPfMW
KSnYxyQUwnd/3nyEqNhKRnpw/vFUewYwTGxTuV00neOCySeWLiA0z88bD72c7awt
50XH3F1+XeX2Vjz/paMLbWi/dhlBJQVLPZk4NDDtONX/iGRBVfkrtGqJCJvHO1Np
BVBATT7i969Bo/w9MbmEKWpB5WRfhL8dpxRmE0MVa7ewAO2dP+Nh2yKqoepk3hwZ
2xHJ7pdJpDeGInGrZTRCIYdodT30Aiuuvg7Xq3rJ/8E1EX82VGYcCLiLs7Y89D0t
pY0M5zmGBYGWFSXTdRIUhAP1BHaWzJAPKjQoMHYmnVKwXVqUSjN/u/9z3km+NN18
Je48PkKZCRfDAfSCDXl6xeeA4iiVhZFATONLYMiwZAabe02AqxCpxFlc/Q0aZVlW
a+LVJygrB2D5arFu9OcDojd0+lB/SMDUyNVtalS4eQR+dGXVJEYzj/iAgN+a/bCl
1L/wIAjbl3MLGhV4LHTvgh5NJ0svZZHMjxT/Ss90jq8wZRSYd7+/oxLjITfX4s+g
UxQFJ3FJAp9oL67rWnm253Q1v28GxUnKUbw2pO82N1YIAQT3sVeEn+fKeluK51Jm
KivntyjDzafrBeP+jsBawr+k8X7FfaCxNuP9iwmShkC7T+1ZbOQJGfGT1pCMhGYr
660mm8MBO3Q+NV8KkOAV7gu+FIOcDqZ0P0uerdEtmUaPJyGH9T3JQDYAenzwcsph
Wzy3scTQtGQnS8HWE7ENMLERtRUDBa1nfNDSJcL5KyPi30aMzsyEgwUSiY7uKE0m
17bQzZrfa+r/vlT1EEZJnKXWE5AZcPS1o13Jt1xzMxvtwmWyHP8jx6wfk2KXLaqr
oHwtcf9Y6aGE/PU9jobVf8Ri64nIczyLAfXadFFjXZj0qfoua1Rmh0ZpKdr6ahYD
e45rzk4yQ+U6y07ubVvNsX7dgkEafEcQdZxExMHyqQ3TuEChTQ3IYccT/jTJgt7q
n4hj3P0S2FJ23xLcMSHK8jlPC0Ucj31Bq1KJgSnZIqTvS8FhKgYH3A/iH0MOsu5n
Wcd6+xixqrIe7HPeUEMyJ4DkhKyAzVTcA7XJZ/Fdc7SIhjHqPN3LAOTNJaeRoWdH
pavMurkmr0BOUIqLf6d985ZX1CtPcvWxLoLPnXI6gyP/NwpLDxsuegcUTaIYPUST
FbmZxNDWuc6AfwWTkYl3zfpxHZmPLxTRsPbPp88ebH6iOFLp1PRMliAjg73OseLf
dIkWkL5KQIfuEbi8ZsanQ7Jo1hEunc4ftPt9xRbpfV0/9JHxwf4XhclrCvQEQimf
67OYzHCtd2tkZK8EL6CdXqDvBd5w3oVz/E9t91Lq43WEPIvTbfqMVztpx+XWPyGl
c7HViEMa0UdQ0lx+5CkRyaCBDWU1XdePKsBB9fUSAVZmjX6RgV0rqkOEXujYeMgA
41OVtvp1wM0lmu2GVslwQ9yy+PKLHytQmQJ4rp/f6SJNTiJy2wFyfTnstixoquh7
5VMhFyTlTT4da6pW4TZ4R00RyUBNrTUtfF+OgrvrmGsX7yZ3g21gIxQPg58eueZG
vbxKeC2c1O5mixh99pIRSgMuvdvuBFIBqMXULezsN7PxCNW/BQWwPWAJD9hbEIu3
bAcz8AodVlahv6cVEnAeBVGaYYSUWqG0LL6enRZ8BdpRotwkqDM6Dkaa34GN2N5a
P+U74kVR+SHUkTHfqGPYUf6jQbo7r2kLJ/RyW8fxTVUInhaQlXDmZZhGviIp5r8X
gB4fW4o8DWc6tKzjrQpPDssZKKIj6t+EjhGa5ccCJbxL7NuIRFfVwZ8kYbs2fk6f
ES+xwhRwHtNx8ekfueMa3N0AhR96Mpd4ixVb5KH6XPSOjf3HXgnDFTcQnV93CrRD
m5MkRAfZwa+4ubzsr4w22LdR0aj7+5ys/CtQdyxfW1fuQmbeyT1oo0NPTbCwp6oE
B/YLc8za9XvCYA/P6hSRbAZJKtwFwwEYUTdmbuQ1a0PmOJh8zwM/ZYpWuDEe/yaw
hmUm7WLu4KVNYTaOm8JLflk0AE/eUNfjY9O7wjXGuA+nPnDuxY4F7RKv2k2XX1B5
2EyqLTMXtEeqDiKpgWXk5zTW2YvidLluSCUy7A0OfwBz0WKszg2O/AcyaWFjuKCD
Z5bigzdNGxNGYCu2oFUdPqKKXRrbu5uIhwpkTb48LK+oWDmd04zV9uCZRMbh2+l/
90vlgEZdMvKZdLuJsVRv9FA16EXNq/adxdBgHYZby8YaOvOZj5/ok49xe6Ucwwsw
OqwAdTx+NCGko11Bwp07Z9Bbhg+o4R8w5KtVQjZMeDbHOH8yICkWI2NigBW9lRsn
OxzFEhU2ROKZpepJtBdrKOvKe+mFX9qX3UksKFuG8byXWEwGftS9jWsfYBsBGvS9
v3aoqBRgN18S//E8lqNvsFusEG0YsShEErKNdfgkOtqsz12rJs1QpugGeDH5DjxC
zG5RsLhSDge23LA5XgCaVlQ4R4vAozzNYJHu6p9Hw4pGJ+bBmQN04qrrxn6j0d3v
Lfapba2ynG5jpQP04kiDH6pEcDAjCHrkBLTLStmXnNF7U5jm0ud2ShVLru50Dayp
qW2GEA1pYkF/BFe1R0hEKjyrLLHw8cHHBMLVINsd0eg0ijHliEsFQ9zsYU1e/wPk
jtFOiyzqeuX66XB7PooYNFG3DOkAYegib0mnsX6wPZPl6HP3sOWT/m7lF9OxZ+m9
xc5RB3+LkU6pBCVkiEBd/ZTZl8cq4HISHFSLcT7UcvPfvLZoucy6NlP/Eyjdyfhh
8t5WEZnG+ySdSOQ7R2sRfJs4LwW9w//yeVIDJ7PxxhKT8mn7dfZ31h23rUSVL7wB
r5JyXev2yJXf18gPh99N6csPXrD6oF25Fprdmm8kzqAsgnFnTv2xq6XDfYZulTH6
AqLNwZUb0WT4n8GTVgqm2mXdeM7wRAxkdDS4jSKsm+tMZhJATGP3sC6VyzB6mxOb
M10sojfYnjAoVU/lbyL0ixtPEr5vvrrRtV6yfVP4N7VQy+HSh4X+XPPbyZ2F1QAF
WKOsinEJD8B9XCOu1n30fpgrSsBIOzN5nv9Oq35OtYxVZWgRCWABPdRqDn8aHVJq
WAjtIcBmj5pxlDcReVan6LeIMCob+ALSqirV1jxde1xnaLPaLsNN24N4vUdincPn
XESZLGQ+em7rrMgoEpErfN91sJurN12k0vqur5IKoJW8CisZlimrKumIKZdhESKb
86bVSZDgds3sfVA8gudiKGGugmckdnpUH5TQtv+5hTV+1CqwFKdaWJ1AQmX1fgfK
+xMCj43A9XU0n3WsD+kfCc4bKJXo7i0drlg2IOi6Rew0EmB/mfcxYINt802f1BKB
+tC3SAcTWBwAfvaAMqjZLK6QJjQPYgzD4W009+urJGa2Edd24qTuGfnjpl0LlObK
sRCDpU81VhX+nrypmoZ0it/iutF8+NxdvnAX6YcEDyyDNWdhwjFn7ibgk0rhr0bB
duMTnjHL7AivSMHVMjLCG2ZuK44CMheN3xMyye1JeBArmWeKD0Whogji1nOBaVgt
fCPor/193uN2TW0Z3GURMn0l/SftoqR8ZwQRnBTKzr465aw/EIL+v21ogPmYO+++
vbMxqIr3ZDWtliQUo+s10CtfttbC4F3X8eYk9HcSBc5lfOMe4Bz/aoahuDBM2KF0
hzPh2pHDqOn3T0WgOLmecC9pneyKyrmERFBWLYEJqQ6UjknitEnApSpkD4c678A0
aHuL/nGSVagK+o98p7PNqm4GiFTKvq26d+Th2QRM/V1dqbUAC5TAiyou+eJPJXA9
CNWNT5krQhVSxxhef3/B+/SjUvbTOyoSqkLovY8Tlerb0NzpyJpY/Lb7tItRFkiC
/v1dwC4tKCJxvm09rLhgPkcwZiW644O4R54R0E8Xh6/Pu737y7mthu26kS2vJFFg
i6y8FIRSW2ILpMc0qdwS7TJJcZ/MMyYWGNSQN2b2Eiqe0WWPqLDOx3UjJTnzCCBB
fxcXW/sKGnRCD2Nxt+19eMCP+5xB1YAyPTpZGrOLosYlBs1q0BjkZxbzKUhM5SNJ
495ef3yabV0727me8V7nKLhdhzCT7srf1MFzxkJbYr2q5ap5/bXQBLFjq4StLjac
nhW5Ayar5oL2SILIiM+M0yvC8hrrpZvE4sJPmEyNySHH2DurN/1RwZQyfjY0S4zy
mVZ2edmXXXJoMbluyk17FJsUd9T+UumKkKRDS/8yMt96q9ML1cvex4veo8g0QZXS
2tQpYr3J3+YeWh+GcjO+JZo9rsYB9zMH5nh0wUplNB0wOdDT8CPN61ImypHR4ACt
FXeOQ3faDmCNWtBnElUyfoSh51dqQqIXVb+nmX85w8JgLeU6+LEg+1G9JgYmV8px
IEKbwU8+ZExSgKEikb53pG5hPSwJnsh1DxAESUsBjcavnDCH6cNUA86eoSi3KAHV
gZMpI0SXQLHUIX8N14BaeWcB4KYJBv12hlKCQ86hGyQHeO3gMMppx8lCjs3VNnXK
3h15Id6CGLp5Wi9uIGozlg156NvyQDCJ0M8xXRFfQEvS14G4iYH53E+kvnkdoGZ3
sHzqhyzDYuCkDYsBr5vdXOjr1b1pBjOwdP08mA89PpK97RypsD1N+baLHbN8DTw+
pShENfh6/sLGc006yrJAK+2nqy+UbpEs9guifA5OJWYJkeJvV72MDIt2o82w0YDS
PFc62AJQovRvhdgEbWXaoOEgwOj9gkN4tLvJ/xrOrnycWhZKmwnlzUj/T9Z6zD6e
qecNcpoLAupsd+JetUHumpwP2TWYHQuL4fTA8QhaJxjVaZBnJhqH9j+cmw11Yl4f
kc7q6zWlrG1FCGxzxAHJoBv6Unhhi+BbHaUSFRxuVFE/zggNGRYQn65TJ8uVld9G
1rgjw/tcKdJwBG1+IUHWs7SDj3b2uc9Zxd2XAoePN6hRJIB0kdnlM7/9BB2d5Flq
uw94ZQ2gAZ+DoPUqKCsNackoD72Tcz+HEm6YxxNOClt6iH+h8aXDfDDOReOKzW0D
1Zj0MOwWZk4zp7Mkibo8Zm/f+fFZMIV1YSNoTbwhTPxEbiW29oQR0g28jnYlDWxI
t4BOy3e+biXMx7WThW8mOgNu9dhnhwDC4OIE0hLNO+AkmV+qt6qQpvp0BEwkt/OB
306ivBGbYmR/rjoNJqpi0E8K/FatxHiN7GwftMDQ5Z/ejmwrEnmRSSg+iDOhlzcm
oHp/m0N9omqGMmE1kisWo2cRgPBmtowgfcfJL2+exfFlU/atxX1/DfrixX1swtSK
TvMVUQA0m9mBFAn0QK4aFHUsbEmh5NHjxr28NJdf5BBWoT2aCXiHcV92YgVemD/7
5jD84jh6ZQva97NMOFzY0sehgDifNXdnO4xc3U/2QJ/On+a1Fb2EbiW2VHPxmimN
8c1OS/Z9WgAZ9aNyH37nfBSbuoZzRvYwPe8FW2nzFYPDGWkBpGcvF8Qbywsanax1
i/h7KDsAzY2rCqa6KpVmx4hAWonQm84rY00Gz91DwrABjkzp07GbKER3ohjAa5Cn
av6OU24tYaxSesGLXsXQ9jRXnWNb5TT06i7qW8g9mFGsNcHlOJzKHo0MOTlae+L6
9U7IKLHsQIelppqopUs27JjkXLuvC/CAG1CYGuDyenCgJwQ09FEyh8rZ2KaqAtBC
mUXNzgJR0Iss2RybS304VYMhwntka/p7uWEVDqNIAAPQT5Qln49CC71vSzx6r1BH
mOogaklAy+HfejkEfvpt9pGjSGyVVxyAdfLHiwfGQ5+ts9IvJCltd6r+FCEhvC8n
194BmaCUDv3aM3f5McM3cQVcBqhZ9fP4vtq/BEKIeJG0sww0aV7WKShi047OaafS
9Hx7Mjl3jMEI+LqHfpTwAI+tMfNK2X84p5JmPQSEBPdBkVuIG7N1H832P8lV3Wep
B8bW4hdCa2FFhm3WGzoLMJxun1fB+TCnkoLgz4JP9Eel2m0zPx09wWnHUICC+m6W
/r9mNvsP40abfICcM9qqbWCAbh0zqnSAvvrMLV5hcwzKl8h1mhRRrzlxY0f+Ky3y
bQVo4OE/hHL6BWQYU4PG/6sU10GkmXk/dglDGIakEkSuRJHk10JjfK+65/ggOFz7
STMNEwUOi4QzGjpGalY6YVRPsJvpxky9tcaRFj/NgGay9RYjguSjb+5T2JVWfCum
GUQaVW5GH/FygrjaU7S2cFmUf/4U9ahForluCQCNGhgyf01GXHEf0FOJuBbSlm55
/tI6WGpqNkF/qx/td+nmTZin6XJ+AEd5lXxjqsPFvau92QeksVILbN7REWDuzVYQ
pI4JQlbhUQf5HUYjzrEW6ymaQ6rkIuZLiI22rUelBFWWn6O5XFd3hvjcsw0K3YV7
Pp2Obn/1H0g+LOV0BgEMagRXvMlIB5ZauOrEsMP0zBLiJfPy16y9euhZe9lVI4Hp
yvAbH8yazSOMEd5FYwxwUfbltnn5iB/QVqiPU1Rxg0oD44d9jtJ7lG4HIizlOAAO
p5jfAp0mfOxNsRNOHyfG4JMys0nYeOZ7ixX/DTxq+Gyt/0lPGRupovB8uo5ekQCa
PpVBa5YQSKq1+DaD1jHbNx+lclQkJOMbnLC61KaP8/MxNF+i4b4KDpoMDa9JfoA+
fulOQBLno+skf7GIuXHRXai9dxAIQTpr00BrSqS0JLqlkIRDsWEn9p71Te+9f+jX
0p3SWcD8zWStjChU+NW7UnO/7j/nJwDwZLcMMB5ggpVavTqv/xVzGGga4pzL6T/i
ENfjSxcZMJNUWAIMj8bhdYU3iETX/D+F90qCKAcv5YYYKnqSloEUP7KurxrUUVwt
3iYpAbNX2F1iItzGBUOTn46wQPUouJbmVPejJJGNK8xuHdBGvp2ITeN8cj8YLJJ6
FQ/BtLkOGxZz02oLtuMF2yzkXKR9E2dyD73EmziWegb+vSj0I1b2XkCkKXttH9pS
oYZ1DWtyIaFSvip5UxWwdYdRvd8COX+jLqgg2PT58fWSIlvYUpxTI8I7yuD6eK6Z
uf1cv90vvDklwakQZsKoH2141AryM0A7PpwNuO1j9evdoPVBvcS2iKgOmMDtUwQ9
kQJwAzUJqfyizUlKYFRt53vS0aJQRmaJFddU1KOHsKytl4/ChnNJv49f+ducc8fm
h0AvTAT6q5aFgj770KEj1QE4K039vdlKh9XSvrHhbZ0mOhLqAwMvalXw8BQmjAgO
/xaIsqm8LIIP+h9LXxgxnfDosIJk1+eyJrCrqovqGoFQIA5fOIH1AUcohym8sDS8
On5A8f4NCgdTUxrNPO2h53qJ7e+7gXhHB+EaTY3r6hF5iR0GtFs2lIJlmL3UnNhK
DauNeMqwAZj5qFVEZDR6at6zOGu67WKNl0QmjZtD02foSTb5GXeetT/6Ixz3E08m
Rl8iUwgPc+Y9lG/FjHT1CdCn4WYxcBlEepV8qYMN5i2TEf4KfP0ggfqAkdstJSCR
kpK9Pnhg0U/vktlRgQXVTvoaW6OHGs/9uS+rfNUITiNC70xQlvm/jPyCf1HVHh33
NMC7b5Q6pOwItEe3penav1ngRLaV+PFF9zg6D35BoVWAiG3ALYadeHntBj5TaHLb
BV3FLFamPOdmVJ3Ag/B9f9BbyyVi4Fd+oetxqY4LjHRKMYNmNmf+XspEJFkL1VtT
6DecKQNXgTzbijWM4ArSUMvNdsMYo8qQK8VFixU1xGaIpHD75XVnHkHhfQKsLsiE
hzJa09nBNmh+9I/ewJqXQJ4jBMY5lcbim5VHCT4VB2R+AcwfijB//9bHxAzBRO5r
yRx8XJpVX9vNclfSWaM62xxWHPV6qOrUQrN6J+zZ/ug+VxJ+pXdo8hoR9selmf0e
J88VXzP2SrfQa+i3qi3jnE/zAkAdd9qEq5uniGClM3/blSj3zQYUvkzxvxWQ9vR3
aKe0EVFaegNJJ/nXNzvQXwU+7xAidCUoIXSLOv1rGESSuXHJpSUKSs/ci/wiNsDC
eY3j+Capvqj12Ee4SpHmKLVcXq7DlSnSIRVWUn3xYin+XYNVaB5YRUDQ630fWOnf
jnICKnQybBeXCr+Hfde+rIK5iYwoReQZbCJ013B/KBbAHE46t4xQ05CdC79CGTCo
HKfXOwr/a1cO+GSdXewFKbUFXkMJLPS2aCLXj7jp4PgjoZ8pNPNrfnu5WCt0fnSx
uosHdjD9Xi4/KJ+cEdoa+oUTqekDVnE7Vgcui8RqJX8fJo2XG67OqLGItVPzBNnH
sBDuF8hoyP5F7uwHkorSiXOJszaFw6cOlkzLr/p8GYsitUxKsCud8XiCUsMQz8n1
hfHB1ckc+4UO2k4UrnVwwMMCEfbP2zz6qNLOhTl+Xh1dSy2ZyBnkmLlgw7xNKREp
EHVc6dBL99Ynf6/q+pzdC+q3BUQPEu3zyEBp5AORnJinevY9u7qwEsvzHZ6sBkFj
+7x67LufsK6153Bu8NiwvHi2Zd9iGuSZQBxOuA6O+3DT8Dx93WzxNoAlPT6uOVM2
2nBgVhrXXQPTVwaGaud/d+pxcNsYg6Bbo6hc1oNsgsJ/TPo0YS97qAY9tm6YhT/5
1IZKLheZ1SJlV/WDIBEYK40TPfOcwUiZbMc+d0Z7lxhFuN7PSsQHqyw0sAGT3GJJ
eTX7wFeQ2eyEBkNjt0X8zmRChBqzZjuxzES3tVdfcjK8JD215JortWvoWmaMwm9F
+M37qrhZxWJqesIELda6xCaKuwB8oQrnPMHBrX7ezimefwvA9qCnYhKtRSV+u9UD
g5RwGcIK3whd21v5CWBkD3wqS5Rw9XaWLseHFW0Knr5iqNg79v+hImEmTElIH2dj
4kAiL8LPKHOSrB7aYzu0LCvx2zOD/e6mffmsNTaXwYHET+qR8964rwsv5WUz6Wp3
u98SjaDx5yD4hUV5PDyMUtS/92LwNy7T6MZS88W64W17gKW/Iv5Hox7IwQo5ICf9
iG1hIifPdZ0QGGNtscOyFkKsGJxzq7h3vKWBXG3aAw2hm0htMiTkYZiCfgEAfNMu
s4HkB02d3iwe9Qv4Da5wqW+FIi5J7dsLiuvxNg9vsnDnwfRyck+XChwX0Uis4rP/
GLLLqkPt+ieDasnigukQvaup4kwVpGf7E+ktoiYhiX1XP+eb/9JrDJGu4xc1RmyL
+LUy87mUWaNJYeEP3oRf8ZCXYZGCP6eQ7jZ74RfPi6O03b6WXBh/uasKiL8A3JDU
tbl6+RTMbMMpMyK22P4YW3iPqXsEa/niWAcd3M9t8JlyMbXoPsXdg41mmIPJGoaU
O3Qg/ZeEJrfi6MxfkwMxk91zAN0tZ8oh7AzqMfm3/WpawKjX2sRTAhg20lcxJYB9
6mRlP3fUsHbWgNyCVqyEWibBKVDQlm8TZL7NxPZnlhVEYbg0cCKHJuMvyjdGO0ER
icMWRwL6ahaKjB4mSHbqeRvU3nR2CSH+174/5zHcyBpLp0mV/fHRJHjGMzqoRkvU
EZDlbqUqYH4dusq//sXLyL2p4T+u6T6/v5mOxZxavCSPrvwIupb6JvRJPG59Gbcy
p4j4fi/dhvz2qIieBHm17Tyj60Dk66vwd+cKZU88Y+hOEihQmU0lOh/Gvt1GqI8l
QHPQUWxUOUIHZcl2nU03eWXitzCvtC9p0FRiELAXUwXh4cMwiwe47+gaZgn/EB8H
Hj06xEifA9XoA9JbDuw5umy8prhNekgJGW0HXrrJ+Q3AWs/rVOkz04dT5Iqf1rJk
oJp134h+v76i4y4OdfJ8ZRhbP3/by5Ipxr0KZX2hLTQ9qADszcHF5SUDnNqM1hjF
3Kl7SWcND1KMRfRmfMbSilNYrDmb603tXmWAD4SiNhbpD1G2KnZe0zXmSqS1j3be
nUj9XX4VjSfNp6a2jGF4OyupaU4/5HTmnjgaZeHMZL6Db0/poWZDRptnsY/fskY8
zyVgtMRCoMrm/0lK/TZ40OwNoLMyJ6Mo9UgTRnJ2Byc9VDVOp+pEp3XcR1cMUtTm
Na17idy6qr7wphnt3TitP3zfSf6433Tm25AZzCqujlM/nwttSz9PpCUHIgLzxdfL
UYcLAoSsPdPbDZFt9R2m7jQZ41dTGpFNv+M4K/Xa9W/PyQutTZH3oHPgr7yghbJP
5GlSbcKJQdllDT7GQFSTpf4+NVI5sq2Li8fWJcubxvxzZ83RXylx90QleYUiiYkN
luz5hmLcAraJunE2jFlMgY+540mFXYIo8l1DwjrJr2A03xF0XlnAkLeyXPDlYzW6
/SKSe6k/lfa9hVQgwzbBDxI95DOcmRWWmZeP/LR2ZDe0n/dzAEY+C0ITA9oGkoh6
poy4d+xIfFHmzZCC8rM69m/1gFjRks86W9isRxD0THN9Lv8OXwxD/UV9KNlfNuDt
Pl3wCLwyc4V2VB3SJ87zaT69dXstSALzLp3+BmgR78Ko241iAuUEAo4D/4mxyzlE
otHVuoRPR0i739XdO2XYIY4L5mr5os85eiVdlcKp0lbM6ccEsw6U8yXf04IG6tMI
ZjtW/9Xi381zxT6alK3lvXNfxwawfEd/kVHUAtqmIgOC5w7Ko1DO8Yb5jJrg5s/s
upxBo584outVInG5Dq1dBqdNRg3Mjcuj2/mACDGZ/s/KjULhnzkLaDmN6pta0u8r
f1tJhEDQCYJG8xnZBWnnn5UDtO5oPXR14uRHrTbBFWkSyLigonl/TNTAJHloM12t
tImz4zfB+Ezfw2HtnfOJjhHnebEiHYDtu/0AfkQGbp4LniGrtwrNju9jbBqLyLln
c5uObQiwDlgl7s6sMN2AARXkp3vrjtLWbl7KGFNVrUNh4aiG1q95xRDUFsRtMzLd
hm+I359j4+P8hlPtHd5x89sECa/3mvljt6M1/1PSE6ishvbm0+2kASza7adwkOhT
NBRSgswWIVtBqQiDIF1Rtua6SQYQIvNBAZhDC3F3yqZaYnwjAONQ24WupY3I599h
T3kC4BEO5iNFCnsJ4reh06GP5HChdFq7eCc39t/sBG82XhQrUlf2DAA3HpR4LXq6
wUp45tKC2oUmRi/4OMb43jowR+ZLhoRLX1uTYswmzaNiPO+/dciRfLVNQrR/ca9f
ZXq3B58GKcmJvuLUJQyCJm11PvR6YklBqL/OeqITa5Uaf2cKf3HdskjlUmD7b/Vr
JKL704ahjNdj/GJHfv/kmF0w87JqLI/1+2Y82lESCzg+/FiHvW/wpw4RzDCVyQRL
QScHNIl982u2Ask3wPR7ftXaszRb9f9kCYA0yvwhNVl9Lz2XD0TF4y/EiQNPehnb
+sELbM5kOZwB30evHzWKYf0sEUjWFjPgCp/PkI6WJbIa0o1M3/wmbJArFWPcDoqi
BWeaiGi05DJyHRn0CxZZMM+3QHrhuTiEaXXWB8VznX4unopzMGNeX/cwI4HQQDiR
HVGg9DabpqJJaEh/lq/W8uzXVUAS86DCaJmr6ctbCcMnKec3H8LUwEuXJDo+ghIM
WBhT0Y+V8kP75hVoHDpOBvVVGlsMphB5e9W/xqsB4U5H62tIAOLDipcI7nHQJc3O
p09H+0RoQf4lWF0tZrxIeCMe5UNyMWeFXU1FQPjnTgDWJelXMUR7NisxdXRFS7j9
XaPWwG/x0+St5ZE6vC4agkQsko2zpwGJ0qeyCnwudlNfIKt/+J3z7YX2zLpHKXno
uZoo/KO8tmCuRAv9sRmSCaT5SgpNji1M+LsGcp94K0Ysh+cjj7TEm7ul0xAulMBM
Lj1czuhHvr7PWU5/v6F6wEOoV1gR4TFmte+xrzr46Ffqr5JAx5EHxdwbZntvATle
Icyg3A8eyPiTprNwO2VuMJC3aIJWJBDEOB+9yQAYUHEOPL/tyFMBPkY0fESUy2eS
rj5+CUXRd2H0zQnvJ42q2nTXJeGwRS8UWH1NKDR2IP+e0r6UhDYIJ+KrX/CAdOhZ
5Abxn90P99rnsYWYyBk0A+6Q067CdAXm6Vo/pEVDDew3i+58R8A6Vhx/H4CfnM/8
o1sL/hAOvwsiXQjkVfzTbBUrVrpVq3OTPY0exifkWjkpE5LcUv1P311dPPDBu7M8
+Dlfr9kszktxhpQTwYWnc2YtzlWCKUarR7SUMz6RhrAm4vFldV2bBamVfDlc5vni
hUC7qwsc9jOPmdp7Sus7tqemSKJ0zlZio9aM+lZ5QyYVyLBQuwvrWrj9jQ5vTWG7
rMEeuBM5PR1PYh38YdLVRUSoeW/gQwCSh4Ovya08Ep72qxGzgoOW8l/MIUE3J7lf
boLJSnhKreREE6Yi2mTXMoYRCVDZ3Bmn+dipE0DIRRKnpOl+RV9xdCA03GJehlyt
AHmWEDGdlrdoELSV1211I+hdJG5NrXoPd2r+7Nkd0diwzk3S0PyTxFYpO+Yp9apS
MRRnM1zOsJf3SmhIO61Rp4EfuFTylTblgstZ/V9ynvvH224h4ypgweVTdQMaYpVX
3Y2US/AoeEPP1SBubVNxi3c3i5QJShO4MeaKRBRbOBG5WNdoJkUX9+RKhP3EQaur
KtxxNcKRGa96QFyO93E4258e/fONa8BYCerX39n4VMlecob+qLgJskA/rvFiAIQz
xpjqoVm6w3e3b0jGaJgKxtuBxI3GX065c3aE0ChkNxMiyvub7mWr0Dtsi5rL04ua
vWCwelYbdFBS5Ky66zQWqATT/dH9iYF7+L46/uB71amsyE+ULZUi0SeaHkIucsLk
HDW27uj0v66CpgZjgz5IkuJ3h+1UOP6zQ1fmXd/zGf3KTGUNuPoBBoKHVKBRY9oB
BO+g+nbqRs5M3ABM1URxPRU7IfFXBgZEbr6R5p9sZgn+KNq9V1CWmLWs/sNRTloP
7Pnjcjpd5eySiDmXy9+lTKI+N2apqunlLD+8XwXFA9/EKC1evBJg4z2fBSOz4mAQ
xPaJSvH/PUjAPuR0VM0dlN4A23HzqKhXnOE8bicFcbFyVsrC+mbM7+mQ18ttjapz
HhZc/1ERqEBzPQVzVCtV0ldb0X29DpAZ+HGRzFGLT5oTKZB+SAkYqOicW2B3Ph42
J4Vhw0uYJKGfgGTqzovpWPjCJAtsItVUxUmq3vI8aQRV2JowbHbyu8eZmh47fjAx
+OQMU70xTR7AG/4fMsXayvsTlScnzTXp/UBwucWv78nHS1+V3mPOgiy3n7oqrzar
rJRo8W6XgzCvgwsgb9NO0wU/xg7EbQFK0iCqx2WXN5sI5YLWU2eJ1YzDiZ6BqglI
5/2i6A2C+gUdmG+r8VhIX9LJ7YXb3Y66jpdKAxV/KKbSpUeMgNiuxISN32Bn4VMZ
s6G1dc6D7X6aqK+O851WT1h7NedQVxkZkPchLHh3eM5x/3WQu6WF376c0noWuOSK
Kwzo3F4axEXiJUW1o9lAK31RJrtt+wX7zE+8RJGA1FDYHIY7kvaA0uqL89+qS2zR
8HaN/iPGiMf1vJC/HgeQACmwYzixsAU8WHha0edC6yZRJqcaJa2TlBlbOI3d6ojx
FxqJi5eyL7qbHJTho/ztpIm7yEW7dBzRHSjXt4IVCg4aPu8rhGDVAa1bQ0KATDbz
XEi37tKAE1SF9rVxX1aAC4/3GKWfe+1SN0pqzGlnJ2671ZxT2wGtBom0xIzp5B1W
M3KL0kWxEg/F7ep3pAHezdxaviGuCt65A8h9sO07KZJ74PlmAkzWSWGTX3sMUUAj
8wOHXNsIhPBled5PKfoQKa+tZfdacieyx7moq/lIQf9Xw69gSeDWPYngljMAA/H5
6YxPF3AimCAWrMyDwDi2lWie72hZ+gcOO4wWIa82pOR87SN/I3St3fCPL5LAsvru
uESunyQeHw3QP5BPoKiHJuTGLu+SkDRyeZdrSksWSVsUMU9dGan9AL0B/afzeXe1
KlqvwzRFaSlSHBWjgkQjunu8E8TvBzPnAWEoMHlh0Ebj+vwfvCfXw7CaizSvtNaq
GazFGamWdqm5go88lVd+0+dg29W4NGvhP0SN5yO6MUQXuocU9wJzOoNtJoigXqb9
Fcm5cdwMdXiWfhP2KODdhcOdqRYykgq1mVpoTR1g0HcqiDH9lo5z06oB8+L/LENS
XwvZRUEnvGwmUEKgQV64r16XDuMBthiQ6bETwM+dqPhm9VilA5wr1qyQm9744iJI
YKJywwK7U0IIhvXtRUEa7vupv222zx8ZWAcnHG9lnf9cF+o/gU6EUVXZkpd6MSFW
GDPcagMtuuh8EDe09vUm4lH2NwWpcLnAbbILkrc37fTidN0M847twh5hMsX4iaKp
LwIoCG/Ek+fWOGS+swVJ3gNhMcK6Hl7laCrE3M/RjJQ6WHGB+FkiP7sYzjzXt1v7
zHklxOlYxM1C4Xf0tMvwM/Zuwa0JqsofWVxR9ryleNKTUB2L7th10yRO8CEHfq9+
5Ghvds2gga2ciT7+/A8GRgAYe2ocabvVBrx78GCp+9ct181nTTy4XRbEDrwvZOMB
dKKdx+lC3kAngRcz0Jw3s2/VS/oSolsoL1rjozpsUxysG7d0V4KAd5Mm6rFVSqpw
DFpRaqG7pvCSyGB6Idf8g5gj5yBwx/Oxn2mlwEYluB6esg+p5xDOWOYnPEPuMxBH
i7Z2MCigJlBjbD8Wa5eDyn3sahF4wBgUhpuJO4S1gVWY8p1XbOy12g3L+HTtl3yq
IhWSsJTVhkDEHyV4HCTuTbigYudNjZ0KI478jaf1u4NVqXexSNOG5U6B0aYGfAv+
asQ8kkwnv43F/iOaIOhHl9hXaowxnnkmsYG4SHKBa6qX5ou8rIo34A3Xnknekoeq
mPz9BYLhsx4aj7pZSaKq8Xi75wZ7HYK/4LTCMnNinr45FGcCxoMGGoPxprpc7M3k
dNkKdIBPiYUU459eolPOBGuY5Ka0Bqe+WPgIogscnlrMOQaHfLUJ5cGY5IzuuSL5
z6/VpoIG0JY/tUTb7V7SANSVl3bBREk2SQRdIzIwCvVX5ghbcTbc/SB6sunKx3om
AWOMW0eK7xGdgN6JPKyGJ3m1uvWiP+k6XkMdouGJqwdikYQAPj0U2M4StLBt6K3h
Gpwx+ryhz3+6/DXaHSNMbe+Nv6I3qHGhg/uRfPVQmg45JUKLQe87dtB07C1mWfvo
P/OmorJExOyqoV6j8r4Gs4PfMcIwDfQVVddyCj+7tOfj+wcwfnKZjxkYMASZRnje
k6uyO0YtvhrTzPm4bzh1rSYy1Q7bzTDs89gqXcf7PQygsbsN9er+8p+HvGhD+ogg
YcKo7wquamzTfgSWf2Fas4Bu5xY+5+JQG192ubJgi0CaJ7uFkeys82dPpCiVWN7n
ffAEKuoVbr3GN2QTcSKr9FOEmu5pMtP4Gf/ChIJMjBsGKT4jlDtDcUfYRMqMSzMg
R+WgfRgEsVKRpKi56ZoWPLlSTdQVH3bzI7gLPFgE+y3JMZnxsK7Na5GKblsqInJW
gc+EQp61FZzo/G9Lx4L0PcGBh14P1kgwjvOToJNz3Vx9AoGYPdA1LRKb4rNr681R
agBTE6pXhdfEQkf2YRVqJww0zbjRbWsQg8I3PSVAJ0ZUovxPkY39tnp7bCujeQdU
8T1fex9BDviY5Dv/vDR7U8MD+zfYulBSbZDVxhiqYWlGUwpExg1OdTYXoF8jII0k
ZXFln6EkgwesGmGIXzYH2/9yUyb5neLlDwedZAa4TxfpUq6eMqkyuXzD42N5Y/ky
lcBrAVCOsbsGgLgkowN97FdGz2I4GFjOk2WJZZ32DBTg8YhxpEY7xJWMjtiTxUwU
Iw9Lj2I/6VxDzMRiEid7qZ08yNS9QQodKmg6UzX0hZNYPa4oWx2gZn579q7rAq84
cUpqmr+iZtdgIKrsaZGkr8UEnIedxGTQ8nquwAUvE5/e7lkb9TWFxi+Cu8yHGOhX
eZkK7yPlckPjWL8lud4NEizYHTJL+MNSYsvPpYxUBXUR/rE7Frc3+1WklXnDkqAp
z3sNKRpL4db9MXY3SXeMXbd4CuMuKZ4GcRYymMa+DeJoHJJ534dBbfMI/YoOQoH6
bghOaB4uPv3TOAX1BemMbG7UpIQec68fZinptOkkCmq1q1Gbf2iiRKRUBrRqPfpA
VW3B+1NI7IVkx0Bb8+qLaelTayjtfHA3MLoxZizqi2BcCUiryTLT+yUaBKUTKdmK
F4o3hWhhRn0XFrwfBHmEhcyyR6rk9jjMr+q7iLihnOHSc4kiKTMAwTAi3+y9ix7M
BrG21vWJHzMLKQib9E4ERzO/rE9pdVemrYl7fsaytwYaAaFR+8wUc2OQ+IWHkTNo
KwNq9e6xTXw0UKQt0+9YkXxQdvhSJCZMwdlG3sDsBUkx1w5EvAGAhTpIVWZBAJsX
aFESTMYTGbXQI2u9frY5DyJd5042Q+v88sGgIX8J+rORB5F95zVd4avcldGQ0QbH
TDRU/vgRSfPzdQq3zu1Q3nk7JnuiN0zgW8HYfNpHDC/JjDlhlzej/pn3uKoRVzEZ
iRfgQHaBiWn1nwU0dXHye3ue1cc2DbuF7wPnGEGb/wY2xoeD6ZdsBguInH4MK0fa
6oAJKMWYW/2pDCGI+BFoEnTX9f3M0DyB/pclvfQ9DQdGNjp85z3aVt9r42OnzfaQ
AYvdzKacoZ0/DMOVTJXXkWyYvNBBbXMS/RcWi4y+BAJQLmckr02c44EwuWKbFUC7
qvB5Y/3Z8eVWx+sFQ5OZNFoVdOoH9kGRPNEBrKLlQo8elQ3L+qDkxLy0m7PQ7ca3
UNlyDagCDAmhd1qdCX5x78ztXWSX+JUXTj6lv+QG4xyBCV/JiA6qkGDiIUzFaCC6
NwKZDgkUbLmIO4y8g+BkiFgtMy9lG0PRnT07N3dUjrnqXmH8yFInwM+stEVB7a5y
ybXpx0d3Yw9QLOCLuAVt3OxoYmUKaO9+f3TJtzL4kWiR45n5vc9vyT5TfnckhYbv
YVDPKfDlYdTRQyVve92rI/8ELjRloYNZPNV+3ZuuIrC2pJfdhApsr50dXWwbZKf0
SdxW6zLjOY83isogulME06AQOQIH2ynUND6dQJ9xXU0CKdr4pGsj3GprrLuLwj0R
SwOl5Y9FVdEODkRg59zqh3ncDlRNLoUaA54p+UGCPybUH4w62HQcVvTlVxdVItPi
yvVNP+wqVnw+X7jxux95NnAILy5tQpQlWOEkIKGGF6p/GN3PsPvZE1kdU11/BKOt
koVfOVAUjj8FXVFj+ilafICESEHqZtr5K1u5CFa0ZAuMf2ibtuy4Bcd6R4RbR6Nb
ozNAY1pDD+Fez1pR0wn1JpmIRaphOKBjUcP/XaRgB8kTVShRMhab2BV+DoWqUEUM
sbiQFvXFLUIWMxthreSgWyKychqnBwUyxQAQso60BHk1R3IfuyciNR96v7W+2di7
JZ5dYgX9Wwl3DlxHD73xE5tzevoRDtvuACBvkFbMMOlkFfU0gL+5qbXEtRWABwhF
g+UgqfSdXD3FlIDVbXAO1JbAj5G6n+lrEDXKo07PA2r6u3qeUindHRFkmocbmnWK
1w7Vb3chlQdRD6hnZ/HK1wCd5oJiznINiwTwcTfIORerNwfOANu4qUoxtvcVXjIP
hNypkyPDxP+/jrKROnVJahcmgqQKzEnaCRILr+OhyTMCjrvEeglVEpLdxfImoFW7
foUFY//aolMIQEGNWe5F2Pc6ICmobpTMqPDhJZ2aW2POzhsaZgJIY/zeACFrFwJU
eiv+GlElQW5J/mEMsfAZu7SYK0WnYL0hCuWOQgyX1bkzMCty2DArdIWnsy86djY2
9JuNJHlk1TZq77dWmh1+Xyi290TMfrHweg5xLZ1xWzFSgE7KPex0JYw5fMu0aFw+
y62aPpTjylLgmFGp55r0GIyClXanKQFQ3G6OMBY+oaaq4+ezJ93czwKf+R7eUQfl
Ov9zlrBpdosyMmeswrTBQlmgmyG21gwvpXcz25e4OGGTzqFPb6VwAVTcBA4RrTIM
mhw4Yp1XrodaSUJzpeXNKCMA9YftUnyw7oucb6v2DxxHXMQcYqTr1U+SmZkNR6g6
o06mwDU3uNq5OFxLC1ie4vVioIlJksG4i2hCzKN9/uj4cMWteh7bFXmmXRAjM1uI
BMJyh1ZT0PTA+EZ0beCKDdh4juj3Tu2hS8fIfnne24iyz06gLaj12iI5qw+Q+AUU
fEEX95SO9HCUSknyRPBlVtyrusigYWZh38Ij4tXe07bcaFpSYlGn42gXY1WBaImr
F6F671k8+8wqCZAb0vWVsRwQ4xb29WayQx3k7MTd9FIhFK/7B8TZpNsROPPGi62/
Sm4EwzXkciQyMGj0ydf98kzillfQzfViL2ySxY0NJxnxeiuVB0lMdTXyT73xwbSd
OTvg61KGFjtMune4T2mmMxZQRQzsQ5fRmQYa6vn1GLP2l7+NudRvv/L+Omuh4MWF
4edATivvso0CiVQwCF9L9BDOrZs5Y8RME32zUlK2LWr+wXjPg0geembai409Kril
YEkc9ilVNna0qy993TniU+B+zVT7Nht7AlxcI+KIWFcFeJsUbIIT06kldQk4wRPa
BkReM2gO5wsswDi/3aqruB9p7hALRr1zOo/paTbx7yRvG7/SdOZqiQeEClcl+GVm
Pqx65TQw2hGJO4MyJSmiS+bIUteMr4I7PZ2/kWH4NKtirhC06tCGCKAZqn/VCH/D
soPaTvU4l7MOUH3oQxwC2tgFSep3YY6h3a6DV0sa1g/qPI34xbmm5Y4hP+gzDzm8
KOm9sD2DC/HyhZ4ocpVr3yKagQL4IT4v2A7ZJbzPX4nTHCIh4vRAo4K+1cixs9rS
Bc2LN02jol75s9l2dJRYhAWa8GzBqN1kiF5gy0n4Wp3de9P2ba6Rf1cZwZtMYDzu
db1VtT/ccXJqlYvz6zdL6aP5VzqHL6wzeMksQvLw4TSG0jvg4IJ21FkgQXyQR7hR
9gpfmzk8TCfJ2RLx76jVPpUzYH9AG42YGUyIbfx36urEUTi5V0FQeyXCWTrhL1JS
Yum+0BtmLy9kTfTqLvpDyWT2I3AwQWA5Uoh/85xfK1iSDLv9Cdzf5/p0nlHgyPAi
MKRHX41xiAMCRUlYOf223jcChFa6Bz3NVhFwhnpM5JNzTMNNgNxIY33pQxg/y198
Es5NnHpazabMC3pPz53BBL/F7kYAgZ12zJTRwMZYskvxu759BSmmHI1ByVY7wkkC
CB/Tazo18umsl1Nuh+Qu2rhp+mMeutE0qxxwV/DySEcYPlrBqYugvr0SfSS8hIiZ
L4D0oVnPKByAEPjxZ0AAsOfoWq5zdZ+TL/Q0L+S6nqUCMhw9C49Y5HD1pY/iAPFK
CRExNrNJHU12S7utJwX2vetE7TIqBt/CHm4QWTQrnBPIKtFqTrYCfp+XnvLXGb9G
rX1YGUKP/M596zznwSxmczBACPXdAl0FQPYm+7ePCoRRYrdNG9jAQ6x3Y6V7Toyy
Z0V+zQLnU0Djb3HZ0nNzPIYhtGu7KiM0k4IZKCFIBN00oG+pB/9gTykHrgzA9kgN
Shj3B8XBsfIrTo7NEJ+RfGhqqwY2qHN9EPa5f+Sh/0PPTUcAPBipmZOpi53GhfTB
g9JkM+IAHKBOyo9qYp+wOoHi7DbyHDrDuDw/9pyCyQIzbxUGCfUJpAkChUMbaAhi
Wj1Vwc53d4vqGlfXYhWbo2dQztzwDHf7qYd1EOKX6fn7XZn2cteoQcLGEfuRI9gI
cX76UVDksAVceAvGE7RACpg4ulo/PhEcPs9oTCDOqkuPfrtt+x4/jb5mKfPLRziO
stAuIMelh7KoS4lT1qRiDpRK84fzE28lGLo/Enb8glVolnwVChCBNz74udadc0sL
FqQah8G6s9p8ZInhEWadDoFiRnv8cnlyZM60LKBYQLiiMbpM4VGdQQfh87EuWFvF
Aq1LJhnuwMzeewQFwfnq48F6egO4j19mgGmhWj8Tw0jF3Vccnhus+J1MzioBUrCp
hFATrMyNsWlV5AJaRfBCR7a2fM7NxXBnXxFn8xGPLC17sEa9OLwChFdj5ypClTPx
G2xKIDqlBlE11jCy7UhLQBncOYf1ET9CTxQGtl/HoOkOlx6cQYWmvgPC5CCigTiT
JxT2xRex9MwZIzF0lgxC9QKsM6sHQSEXf/Ra7x1Y8xgjrTmWmTaRMrdSa6VssuxQ
Go6NAAPRrCEIf0HQf+WANxU6S6Vn3IGvFqeJKqz3mRasJrvDSnLTSiA1K9ndgzkE
UrO6vDCovOaNDhKLlL59x9TDDDN1Il2P7hBnZ129861w7dABvU5hRzptd5ksCVnV
BdftmbmK2Nu4iC90SSlQq2GA/CxNVK0eICnw24zyGkhTXAoz/UQCelBWPlIOX78J
18fyUS4BE2E5vEL+u9pdCeFnI5UprM4NqUjr3eyLKoQsXU4UIT86uw/HUaB4te9t
jxRhfEHUI09T534jeo4wo3R7frvvxeUqeCbR3FizR9DD0P22iULrHW3w9xj3FTQ9
T7L7feIQIj/FE9Vho0S4Ci9OJeSckx6MEL5+866fWuZTwiqwHACRl/3CxGd1Trfp
JidK6K4vq4BNhs/o7Qyphu+R/Hl9J0cq6UeWra0wcCfNKZNn0q9TiWrMX9cGgmkB
jAMtwnF74oteuWMgqYHOYNdOrMJUxryre2YtMpz54cAiM32X5kX6PV0UYnk6Cwr6
HdWssRuvKZRgrXLp8OyhibOG0vkkRTRFYfRMBDoo7itt7G0wWKmEQdWmn8Iwfksc
tc/6mpXnS5KerjXJGD1JrDIQWoYvjjj1+vQkIMqynLRrRSGQavOJU6e9u+u6debs
aT5e5yC5xpVZnP2PssmFm5EBgs1tYFVkUp2NttSWPf8jp0UWg3+JBZ2nnMQqfw/O
Fj/+gKURDRpd4keXue9mh/c1nT6Qn4vYj3DnrHRbSSRuA10tXv17dAalgR4jxV5i
HHzZKjm27bCsHu0IzR1YoQ+5Jz9+Sebu7e7Ru3wx63l9ovoPLOoYcZjcz7qSg6RF
aBj8+i4EUAHbLQs5z69aJtkUGVQzNEk081/le70inyktLWyl0vQ6S4ovJ+VAviXy
l5q8XBRESnHOS2Gf6ytX0ZfzosVKtSPUboYbohWNYN9XYAakimkyYZn1+OMvgb1h
S2s4aOaUfAjAByk7HKkt9DigQBJ85CXEnu1tOOxqxJoQNMXIQInXyFjzh4hVcGYy
UQIHdbncgQzasTTqKfETR8BwYox4zE/XGvQmGNo8PefHgRIHYrA2CWicz2DRvTiv
YfiMNzyojmVgps1d9z+zXDTSc5Rg9cLwiPrrC1O9bd2/y7syvXIQN+QoM64PJkO+
3cuOYZpfYxE/P+m3CkkOip4vSa85CSP2TbKsaKf5DtVz8o+trVEPkWJWyxVMoyip
IK/YW7nw+jV+EcmTx5aodaKrEO/SpFMbByUvn9VFX9NizYsf9aXfbwx0vkKraiGG
67RciEeAqi0j2ZTL8yeEdsgbPC6/9hgqoBRT5kzvmpAgHvdfldI7BUUL3Q8vMq6s
TiBzxXuk0+OBKuqruvNQS9hpzG8XZmahe1cwMCfXgBABVlp9cdzmwA+/e/dLpGWf
2A/7nUAkKXsdnMO1o6d4xKY5WXLBJ21640DqnP5wcCbl0qEUtB74YuYkiShfM0jz
G90fXmQtUenCfisHd0axfj36DrVPNi2XY1fPAbV9jkB1dbeiovNufTm5/huvIA5O
b2IIeih7HyMviyfOoSU9Iskkk7k7k5pCF8e56sCy92YDjOHAjMjr7Kmwlj64eEVe
3gL/Z1YSF0ANgUcuyf4ZQzp58yxDNgFp86semSkNFumdztUKWldBujFBwTfYkLIV
krfhM/DhYO49bJ5Yezk6mIf8AwfNT6Pb8IX/LsqLOox14mDa/dzIC31vu2d5HjQx
aZ1iKwWl+oK0RVWD07AqRrsvW7yHV5KdrfcTTmzL52oTxOQgoC+KZLlIGqn1KRST
n0rzgRZXlqGcuY+pmSfHdJ8Avszfpw1gTt/M8I0+l4ZjDFVqS/hBTdObuaDx7dBB
1nZGt+nL59riqCK/Fnovx8fWyPlwMmwf5AJI9DZhcQc7ME+jh3m7It5tm4CDx0cg
9ix6WJCh19P+JISIcdqhioW67u3u7FOY66fuIIHABxHNySYyyCNjzKHOX34rKWKW
RtIHnOs5a2NKygnXnWWG1RXPHcXbaOwQbz5L4SQg+vb83IW32fMOtroZpw2f+t2s
e8+wcQd/g4CbEx6EbPqxKqjVAPYGXwXXqd2FvUqeKFwl1QCzwYeIwjtQIy9dYz8i
OYfULg4vas5QxoDaKaD7IUhfciYhjGRhQZCsR7lJe2k9e2WCItUTyNJkBIHd6Kmj
pX2X2CKUittjdjNY9dZG3LtEeAhgIlsIpaexUhjUNJWjCAFXn/jbFuZRrXcA3o6w
p2OPoh6OdfYud3GEgribZ7ZokqQL3J3JAVwtpJYu3z996i8dNGi4dcAKTGCwJki6
8rwMBghrhiB9fTCJLfVXSIg2TW5AXzFN5pxqz0RBPVSoCb44qdeeWHhswFI7qgRv
6vBzN7H3/3KeCeG4HJyykcWU+Y5wLgNdtEHss1t0p3RO1pC12W4p1hSnOsfF4647
ianbmG8Ye7/cpnkyZsCncWvP52hSa0ZA2JJyFdyMq+U/mfOiumTxH51/EcqUyGIE
K7/1ls5wbRgJlnbrkdffn33aOCyaoDw+emmpdTnoyXvTRDO8cUNzK548gKjwOSnU
ik10AbWuYXBa49E6bPce/utqRqkkEwtE8zRa7RKpHiS49mOjoKDdG6er5r9MVcxx
fYCLEL5jf6iXRucOOjt+cMphngKpEojE+TMYGm5BnE+LU4iZ4rj0+PC3EvCrbMGy
Y9ky2/oIeoLeEDHDZGsx5yLRwJsh9hIxME3YbRmC71u6uhrdUID8Z2LcTDQXodKS
uZvHg3grX/C30c1X4tXPK1xNp4mruYujEJCRdS1mxnXdrIEdJAapMNn5L7y66inh
ys12WBnfDGlChITRZrrmnefDg+ePHYza6dY81ZPFeVTpQA6/yhu9xzQR2XNJnJsG
1bONHn2l6DpY4qe9W2O8QaGc8c54toZE18F4RXtzXtu/EH646eLpx4uj/FU0fsFm
4ZtrWEeO0CAkwxmbPMvyH9xxlncVLjFFZPkdfqgcKN3uKKX4AwqcEt19IQdmSnYR
7Oxw72LtL1FZGFQT1ryIHjEwHYu5Ajoj14+/rDyh033WknAC6dqrapU7pGbM+Paz
niUlHDD2MlHnsS75a0kmcE/TbmWgfGq3a2LUaTXqeqLkQCIXCT1FEKgYWFDG2npe
0rftO4M70Wme8kHJe3uQK+3p1if5nBIGmCkrf+JuY+n74C1mbIEiAMD18HbBFZNC
pPLNSMCKoAf10AZl5zGbsJEpoTgoygC/QyFa4ShIvXSZcy6IZqbx1cEcGoRV/UhG
ccnmu5tVfozKEZaLuDcsdoV96H+22aWY2NBEdMDoz0122uo/LULeuoGTHpdjD5uL
BgZh9f+lm+9C7wN0AXrslHbS3sjLncV/J68CohmXmP/onZgyLZq0JbcJ/jdUSqgZ
un99Ku6mFp6NGa7JvMG3RNugVFOK/GJlZpHbxqUQ05Mcd3+aF/zBsrbKiw94c+JR
QgRmB8m6kMknG3sWrM3MSccpCgMgY/EyBLFf76OgIh1R3Naf3k9Zi+BvIlHVphxP
okI5JcmlVtxItmUs0oS49wr9gj77uoWDHfga6csWXG0+fAYHceGeXzDkiD9Wk8um
Tm2lYP4Tk3EvD8a5fr7pXUHRDIKzoDT8VY+Eae3Y4EIlSotX93VPWhqSmXc0fm3U
1tqmHVnhfLkxFnNN46gnVmUUe/MPFXuwifA1IqyaH5vQBewce8GL3YW+RPgMmXmv
wrY8FfNtsJu2c45R+5pLA43JqKFqXKVn22GuA4lKuihFpKZzQAuHDtxJphrK/J3I
9EtAntWOoIMHV+Cegwx5Xe/OrqLmpTAOoGAuakNhlfTWeuYwl9Z8brQsJyILuCTY
x+1258GAe2VrSpqLpY0mOwMahH+DXNTdV6wq+/PODDPoNV+nE+PyDUvbnMz0tkRT
Xi8QAuhLmJH1MIA/XCs2oVIAYymufXEu8FSz6I7Id7wR8xb/71pLwbTu983y8C8A
99OkDMO82w1OtwiNM1hUvGBFdx4Huq97zP72O428ih7vzJIJ5t59NEaCUqiu97bx
U4cCTlRkx/LpidlA4NiJMW6o3Yk1zk1K2+4S/cu/jqnP4u0kG/1m4YNtdEXoqG9r
U3axpOZUxAg7Want8dxKYjo5m6n4Ob6xFkFpj1/h0oObLZV90QyMgtkhXNxewKYM
OmvjLY9GukBn5Dt96ULEt61lYPEpLqN/rQO3V2vHnaNLX3uOwDkDVy71TWcEuWIy
wAqZ3B0eZHWW5nToikLnQkfMdTaseAMW3sKCM8X47LMjHNAsWgtQVHYePwx6pwWH
GIotnprbVt1UsmaCpU0n1IgbYBMqqr3RMByZ3YOhSTHuvI9sV22tEPFcpeib+Pt2
IjNv1JE/ZcUie/9PNiiNTIuctxXtYykVcbhEjwa0IvC0+OxZaoqB1wHYY+qoowtG
JSJfvRhY+xZlAA/2Kly4JP1TfHpJOFXe3rtrCqizhjx/AoV9i3P+aLqL9+vdYkb/
TKz/7zDam6MxSoCoFv0ynB9w3T+PU2oMz+kcCmo9ZHEC3nFtSwY1H5rF6lfRJwfA
/wExsLf2qyF1MfeBr77mMMJeSiJbq0f0NzBIjJYo+sDA/v/PiEoGPLyge1PyYAJO
OmYfW/q/IgceHH2gVY04yWfNAFgg6s+Scuwz0497bcuTSJCfOZRrmkSPRz+4NWzx
+ZmGmD07iwlmiQD3O61hHAT3iDBZNQLF42QP5TAIlo0MDOB1LAL7F7s3qrWdsF+o
p1LCCErdRX0r0JZtt7HzdrufKNiZUtP6Wd3KWe1QCEzvfeXir+59mdrKFMp8A8Wt
6XWIQIOlVlhM52ZJmcN1J8xgWT14mdCANYnGLg5VajXwS5zpfPjzIjp319lAPY90
tzn6+h835rIMcUkf3dFK1sTzh4l6HN7UVhREPIL4wNDqga7Vlvar/Mp0uQ9Tk81K
MTTC+J/Q/9wpNmfkwIP6A2unEA3x6+fs1Qt92yNAc+qZzGQJM8B13SnBpQvR6t70
IVYCDztmsM8pTkFvNwTXCfN0RMhI8BSwqt6opQD+arf9mIV8Sks2GKDQvBIdwjKu
b/FEybOFY8nRe2uNEJcnGj2rlli0itqoPlZCxpdC2aNK2HpbZnwJg0AjA5HKHNGQ
AIunMDq+xZU/hdl1csaLEQYSLOnj4WtgC1hUBlehkjMH//I1Qgc1M5FRAL9/HEQ9
TdxB6rJeskblzqkYX+Wto3+QX9txtUhiY5HcAFn61ebBqgsQQD7Z4GxzQI6zNx8g
v084D+s8I0pWnhoFeHHFZ+gqNMHBbCjabjrzgjBnx/8AvSfAlJIpKwAlFhl7aqsS
Zzl/YiosUadjZ2FhGUC1s8D2PEKj/Leg2uLndGVGKGze6bQ7KETBYjJO3SU8PIHh
Dg0LedN9WJXwp0J42Jz9WtGjc/Zuq4AfjVkrC3i5CAn+JmdYnvBlsKvW/+veWzU8
KOFNDpekpmdQjFsd6NlCqrEi2mgsQroS4TUJNnRPa+Z2Oqj8jWCuePotFM0y+5Ua
j6NaAXDqlVsFFNU3Mysf9dQwefCrHyLU9L92g1xYJvIwcpUFsskz3WFU0b41lhmD
pTc6+pPIqWZijCxa+3DW5ntiOS+25Z0joqKtH+EVLmr4kUBJo9upGuZzZfgip0YX
1odJYHgCPSpN/IBjmZa3xxFzvKmiB7zJLLe0ZIrPStYRo3hIlnT7iIUy2D+1tn5X
rCZKZyd+04QVc+KQBFX1+oQ9hqTQYhf/XtnRh+8fISDgHJpd3TfDiW9NkhzEL/x9
SvqdPflJrgC0gCSgHsGUuRYh14typbZ/BTKMNwdvC/Z/OVCuxd5ZpXSTSuuBX1Yt
7oExOxwI+w6EW8A7o7VBoibyeSzhMYdytLsmVc84Ayv7o/Yg5kJJAHp2OpBDizIG
K1KEkA4y3xvHnAaHHHr5sscwKaGa1CBxDY6YIfjkIxlb4SfvfnGycB8z7BnIpFVq
uxU46ITW65nf84ICHcAHGv94Gw8KfSdCIsIPcRofTKeV06c5mod3VbjfGyWgPAWi
fKFYPwOMgCm1hH54GhjD8eCtgsvsYEGrxfnAZRZemPW8zCFR5To6JzBuO3XsPlLZ
aXpNyL85i2tRPc9pJSTLX9qUw+Jo67O9x3+XwjZ9cSZ5R+/+j2uDwMr+nkSnIo/S
HeCTWCmpnpOYfombIAG4G9RRGrh9DXAWlVAX2O7wwRd7NDu26QOzZO6fNRmj2WaQ
sB7JEMLIf+xfnrYw0Ir7Kgspvy7nP9rTTSHa9pJ46WYXGUbjXQDYsCdFZg85VBdn
ldfcH9TGFSZAuOE+Sj9IT88TZr8sIgqWIq137jlIXdNy0ylXxD06tIdYLckH1o5d
A9bw+nystgeOXersDq9kbAS/7XVT+SMRYVFJDSJFh3Od28i5Gl9iafs/3EitOCIT
SX0FU02442zQiqPpeTgcreVceI0ua4lZ9nAkfkkoeqleXwSfwbt+Bo1v8Y7hyd3S
NCt+CyNgl4doiAC1ukAvlrlv7iu2+g9lVXxKqBlFJBNi0xZyfjjC4JpLnyEvKA36
fVY5el4ClXYEdQPXsfACG174FhhBoEUqsjdixEkfcQn2RWpU7p5+wrre2IxEMr4x
2dQe8V421N7iOUCjFkOG6evgFDFSmo3FrBhFoTnAKdOOTVC+Eq5MwkeNvYyaO5nG
bHeAv73DprJuUiFf7AFIpprpA3cR3RyJtwH7kxUhvqcXBjd1O2XGQQPA3o/rLD5T
wxRHStUpY3EuOFWhdf3GTNytHA9TvVxEuEVq1LE3cRMqmCivx/c87jyFZLYPBepd
wTKDhYMxNqmHkuUp7QMNRpt4q87hJPYP3Uosef/JCOsBUyjWCsdKJFoMRbLyRRxd
P3kv8qS9NUssXWKrnLdGB+4+Rss4QSV097lS/AQ4Ri5XGQvdq7AYku69dN6gEb6V
N8qRXLMLIS4a7b4YGxadkCkxWlkPq3Rn8NTgOw+a5Jd14+WTJWdGavW3Kkp7gRPW
Ibg7wysRdIKew8e5mxpl1GTH1Z3AFgN5vFLAw10HwoH4SehAYkwrD+qEEfKM/qqI
bZchxY8dmSSUk/YM2V0rrU7vemkh9qW/SEu98R+09xLuXaX+ZCO+0/K8/y2pSkkG
SXtCKN2o4qUkEq4II4COwtK45LWYTijhrsh9SL7gttpX5T0iv5zNdMj71FRG/nS/
biN/SyZCPfg7Ywdq9kPqRqdoGmN8eaZX5luSMmFupDsu3KudFwoQoSwKoyZGAChl
+wD7Kxr31SH8Hy+D1nuKIv9y6Dl16sr8hdGfi9VxMu6YFdX97tS6rARZtjBDGyrL
uW92tjKSwtlC03gyi0L9YOTqFDI04k0ZBCqn8TJAzEK010fNpmls7jw3FuMnuzVn
uXNR1FKCu8KgrC1tvjfM4im21QzOU4HxwrnMBGmaSgkBruI0HELrcOf+D4L5iald
eDxrvnQO0bd7OUivWGytO6vYq285ELZt3REvfPPqqNxnLjBvcNJLSfx//7HcrB63
m4F3aZwjR/tfpIJPgRI8cOJUgeQVS8/tt9HwJloEwxAiWFO7QqooH8f7ul8uoBDI
MvSqBlKjeafi9dh4Dd0mUlB67eLh6myLiC8RMqPMjAVwzClihx1jVcCT4RxJBzU2
hEWYdiPfuTjnEvFgotMHyGBM5u2WkOChJkAwSXPxzww29uYSwsIQrsYfAXqiONtL
pkmLmMTQVsniJTdUrwvQuYE7K/QkSmN9JLz4aQm3pNlFrVlXFfKbEjXhJTpd/oaC
MDGuL0dNnTER5oqaYvkCU7J5TpFgdCDc0mRIHiCaPfemR+BQVhezr21mM/YAuNqk
7gVlEZF1X84re/Xhhd+GxbOzUWdmouCOeqIfHUhmsmRVF2znHPA5L10ygRi7cBcb
w1bIdjsVIhDn2AQBSy1YWTVrJUWsyEpk+Zc8C9sbaSgIIu8SZqEZ0u/oQaA5eT4y
dIS0hsbazp3lnmUi1hIiuTrqmfsKZfwI4sTrNYTbahPsLN1Rc9zGKWCUFLUD9CPL
PzjP88rBREzHLKexptvXaOninsPi9GDwsYnUfPI6e5nOeAOET1mM1Vkslfkr0E3Q
zx6Otk1ktMrGD7ZoP5mB8l4zYM6l3Ce/EmBpVrk51hFZ9CAWNoWrS5KqLv8ecvYV
/gC9NR/VgeHjQx05Z0aDm0A2j+qihH7OlR0EO5lvC64WAz+juqwiOhbN9iVZlSQh
2tkxUKaAOWzJDfmOJVweJlwsO6loClYSUiwVYOqC5u15LQXuM4zaVN676VElHp4Z
ZFcuamm94XzWmWRiz6GrP44lNzWLi6qS9LuyWRYaclxsSem1fytzLes3qnVPPF73
B/FWe6/gTNAwC5FWV5cazXJFnBt9v3fF3qIJDNmkjowirFS9s4Zb4gIPf4jfWWOo
kYVFvQ4UkFisasV7HN0INXjPerc4gkevLjxuXWui2jYrd7cfSOPqhfzG8xcFe12z
LbgfFhDFVntfZ3W1S5Lvxz5IyU+VUKyWhgUKopIrpx2zgjdeMhO7OSFc2fT2+8hu
amm5cn+Wm8cnzqGscCQnbLwcWPH6v4KkxsUtBVTjx+esAerKXXp8GhXv4sfergwP
N3y2QhXXQIRUT1vOA3z7DCZaI2F+l1dDJGf/qlpaYvgSIFS45KZ9WB9vLr2MyI3u
gsh7L2zkXY0/JerXouy9jgQdNRCrfOzvSCrs7/DLm4nGfa7zzO1u8PBhv8z/BAQa
tnE9dYJsZ12p/iFxHil31f66ZCkp+L+uPvxq3Px7fo0ivpmF57wiVEqhaVveRKwp
myIns3wPqaKzeZHujNZAmnKpZB1Vvx8+WOeWGIwI/2WMP/cK2sCF+dQjQKg0qf6c
3PeOvzqoI4T2N/htBi+bgKKGgYkzWEIuI1Smy+4P3sIaaKea7ry1givWYx1hy8P1
HZjNtsyTQihL5Dn5Wk6Mnte7nqhUwgwM/wU3hhLn/6xAnNHr7m1bajXxqFy8cpyj
TkmhvbxXUly9g1PIRTwel+tWfD7piYSW4Q+ljIydm9JOAJVNLsXDOb7iA0UHOZe+
jiINr2WFfzZXWsoTeRLFyQ3AGpB7tMbKdYr22RGLvR6uQPktOmQZvVuVxJm+veyV
Z/6HsRmsW/yyxRAZPo1Z9/K4NVMMY9ln1CTtaGVZ0o2HC8YoVjuDvQKm3e9ZNcRR
C5KArn4ZSsSiLxNWRjljwGwslQaAaORgzrRGV0nx8gq91SfCJ9jTD8lW1JLQdGU1
cNBzcGjZr2C/yo2+91rNgs5kp9v+qSKL6DbWtDNuID+i8HIFRPA0lkQsxryVWVE7
BmBG+FLpjynML0tw1JIAYN/3VHwUmmqaUwuOsF5TdbQ38up9ZgDUalaDgzL2lLkp
phkF9YQPduztWQ8OrfSSka8eH02sCvUOi8DV8nREdruQ+pMeZVSdKcnWzRtwb2+U
qel19UUKQDTFr915haIxHXJusnC9onva9PFlt1YTa69eAff9f+NfXx0Kim7rbfOT
jbKDdx+VudKfewa04WtblpAAKU69/2FTZ/D/QZpBvA7Xj4Dk3f2sZ6fKVEiy09Eu
0SQ7enT3laoZQ2+DwSh9RK4S8OXYWHDbxmPjVi52SCyce6Tp42sDaLe+fEfd0b3N
x/qbopGOAfwDs1Y7HFSm/Db0IUOA5jhmjdn/Q2zOK2pBelnspJoO87esxzEmekBy
4Ed87EBu4RCVQcZRGK2xiq549cv/zQjjqxzR8iZEE3z+uj+COJRDXHjI5vg5OY1c
reDigeke+S+jqhm3TDg1KWgH5ZHs7p9A3hUTx3sAcSGQuCNi4fl6FpXCkkzdrJse
TQfHs0wCEYzgbJCYN+DG72dDC/TVT4ATD6ir8lYxlU3vltt0KfvKDK1qT+toGqEt
Z1DceDtXj4OLDUmeAz0VpB5ef3Sq6TKCGXqC3u/d4f/uA2kYMycuWcDSWaOk5DFO
/F667QKTNNL2z7shgjpNOeJ0zMC9p+6SvQxn5X0K0juN7Guo+z77u7DNJqVK9CrL
5eVTwBlCLYGsWajPkCQduBfJ/+tOsOhNK/8KOxcEtiJSPMPP54lnSFKN0oYDMCrc
63IE9BRLBqFGPcpMtV6UgGG3+SdaEGG96NiloRUKWh4iCoUkUSmXtRwO1Y4vRJyV
ZmGUFxVYzFldwZWi+UzIHUjiCv4xXzP1zkzZiXZ5EZid7cLbLZrIYZG2D50TmAEO
sXXNAI2lKuxQpc+Njjzbn/3F0GpmehAo5FXcYqO2H5M7L/pir5wENf8LHTXjFR3P
YlFkcVLXE7k6oB8fnej9rBeQHmYoft8cjTphM742EDhhCLHU40v1y6MXd/pDAcqk
Nr38bNAKxSezzJMPJePTn82/uHHEEX0IEhyYVAqyQIwOSO5Kq3+4iGX5GaVXrZ3e
OM4f890RzTGiVOSbUyItuo0FF7pEpnHX089uW+PAtoqroHeWnvyDEVwiLnVo7lEf
Vn1zl1UiVAltSiz9onnW115v+KWtRZmA+z9R5NqVQO3ScQF2tzqvvNwiJPzG8S+H
8cCngbqustD5GDtytSMiEi2ExhMRR/rm3KMLJ9gd0BzGfuME4iN2dAIZoovwTH1q
NrMu0+L4uRcGCdDZqoQZ7AJfgNEXdqPsb9i5bMDLH67EkdZcy2zxqA5vw4wP3aPu
2NOUlYEe7VSArHxcOPFnF7CP8Ikp46D9QmUz+gu4h4Edwj0fJljvCqyWYFVE9hS8
N6YDD28SZ2bBZSI00XcaLh05itH8Lm93AlySKo/tq6Wd0ZuWd2lwav/6tgGDC3v6
De9lc4ClR/UxHx3DxazYHGUUSyFeiKUC06k3f2oidt0O9dHYxYCh0+CrCqCtaFoO
JfSpjgkUwg6u5TYrc14TIQJlxPwqZNBwITviBliGzhsR94WAE5dj8oTL5Pf7Hk3N
wYKiMBllwS6Nf1DX2JrDrWu83hLsTJjIFxx3CQFmA5qk2jMcNH6DwS0stXNpYyWm
mYPeGY3wdtG41Axr/lmnhCBp+51Dwwzr0scWE6LZhgpz+0FpywaxT5kfyLq/t6WW
VcM70W9l4y1sMzrmbyjIQl/l5EPzqMD/+fL6a7jVVhE8wzmw/827lmfcixmNHfa2
CvenSNHSzMPo2+qnEtGfZaLrTZdXZL115ffjh4jk+3Qlbbv3gNyIx0oRL34QZw2s
/wOgYIfIUQB0wz3NkeIooz1XsJUt/R2+zku3twYITgYMx1t41QRbId25UAA/QEB5
dpE4dzDGBkObll9gzS+7604ZAcg8zo+BRqoq8NJsuJLQJl99XMbn1NRUhhNzZkSE
NR7fAR8gU34/wSLFSSj4yXRu967kcKihldMn1X0GhITlQw+6VRl2RWIBOA6a90Df
p2V1vtPbqsc3CPpTIh9GGW6srAfEegmLiItLQbTHi8j85tZI4Ht//59juEFBzcIj
arV50CcmLFCRk0MI3mab1yRSMCpeSjudtwdDNexIbRLZ/cKjNMjiYu61TAQVFn6Z
VDronLHaBW5nuUfAC8tYzAxz2MOKXReqSuyE3O232NgZQNEtJhzX2wGlgid/zQFj
ZRCLrO6mAjuRnfGIhgwATMGetrhrD2zHxjqFcbLwZ3ljdEB0L8n+75KRljXDTLpw
WIX/njmxkHmUOfr+Nl4OoHVvN8dLVsIdY2ABJHjcsv56bwS2qW8k8arRT+tlutsD
ztowYL50YKC5JxttOcXCCrNOFe9FEgCpsBZuN3qc+F0aj42qTqYi4XGNlR2tTD8r
i/lXF3MZY+RPnyYgbGEgzcrufHZVu10p5Pr7VtoWoyKvt2PBQcpWjpwxdrL4/Plt
tr2W2PmYqIH7IXMJdBha7odtNp1DP3iKNokJae+uXbrv7Pch1N7fveZQ56HI4dEz
NBCVEx3hzYLYyCxNwQs9T5WN6DL1vViZm3ML5io164ensVZNLrvLLC8sRpqC/gVH
BhuyreQXsm6f77UVafaHlCv2npVWWEMAnm31S9cXOBmc9ZkymQAHaaEa7+k+DRgs
kjN4YgyCx/bt0TE0T3OQMfuoYvzGZXVla1gn68Litmxtm2DT1pLiwYMpx5N9Xa8V
JSz94CLcgJ1N1Jr0oP8uUlA3mYPGcME8XqbbDKlG5ByyybVFILhTYz52WvYr04jq
tIeALaGb5TCPZ/GJkDfZzAiAqgEDgNhroSJP5awd9tBSY7yRiUh5Yq1OMfW8S28W
/o58CjN027Y+1fvJyg3TR0Cyi2Q5xq2rx/NgLlU4cPdLEU0NthhvrVz3mF4YTDKz
WRTyi5uWeIdbZwXEvV9QrGlxaKa4sfYMSiGtQC62iy6FXtDeyzBkyTSH2pnNenLS
NbuJnMmRdzQNIEZGJRxS5oDSbV2fvrotlUKC/jxw6/6uWuBInGvKewmcOXKUHxTR
nS6gKa99KfNDIMZ8/vvO1lcQGBBgPvnO+fjK+NldUfB0pbo+/NINntWEGWjQDymW
13ZRRkCegDQqQo0OUIRoHXm4GrmuTOOS9eDMg00MeA6RSmcrBu8e9+1ewFVAcx0h
Ta4IXB4Vdw66zjNH7E8C8IahNXiQS6YNwUsAyJCPu8Yt45PBrRWCj0reTTaQKK8m
2NIUoJxcEe3QoQG2ZU7JkIJ6J4trQ00W26GgaSD51rPFTZrdDVaGfbJiU9bd2muG
dX0lxFebSrbLhpc3xDhCaFu9lHk8aN7grkDcMAZQ8yLNZT5KLzB6vS8IhK3PrYq+
Eyjfnh2B7DpTx/cu4vOINP+bFQUiSPlFW2F5BhHR/JDfIKo9BU1eqI9TVrQ3O1AC
daJPjtk0BCSGdVxKFRBdZsh0kKrO9P+vEwZ1ZeqyIs7TEOwCxRXqb2nmTtvDdj0G
4EgL3Sx/072MDKSmjPSxBFI64OhHchbEe/Yq9d/QkG1Wi2v1KyvuXDMyQvEesRNQ
sIdpAt9mUI9NiFRb+UZRk9yE3sD9Gxmu6K2MVbrpIyrXSig9Y8hrRyKeMsqu13gS
7F5YvUCGI+lQeZvxkdLPszmKmytZc2bRnfd4idHxFsgEScgEIhIQTDdBDNOl5iR5
DgcF55hnwUXOz8Ho+OWmKUKP/QnqfEnnvRYJKGup44afX7fBs0v3ZuiBAcGRxamP
8rUgMoBnNBKPbM1ydlwQ3FVAwZVzZzdM4CRQnNgWbMs3TRZNi0x2ItCU+fPV5foR
7vyEyGCX9lg3yYGecP8XqfkPrW4slehA9vqojKRMuAHUb+FDuNc6E8+j9loeSUj0
ywJRXd44Rc5Pcp7mKzmOVQgp9rQdEeFltqJ04da1Tek236Thp1csupyWU4RUWxp+
vi8btg8PQYTlvmbSfUNOn4zUW8dMEl/jqMUUlJgZBgFU6JU57Z9hnXOKa9qfKsnM
+bOULCcuw/LhnZ1GDbfP57OO8BeY3AyaO3WdWQKU4586a/17twt0F5m9kiXyI/Ti
vHABvwfm9SpjVzpgpBZw7YSQVZYrGJx3ZFjKYUbd71KR9YDfSC6R8z3+ePVn/eIe
ug9hx4rTPJweYmz+m48f6XqwpbMNlIrJjeABc58nrmSgZ5O38T7oYw9pWGHN2Id0
h9qNgyncjnCXxxo++7+kCbn0yO51v+CWqxB8kW0EgMe1NEAb525jUfM48QYHwUAc
vwsbD2inMTAVWZmvxA45aLODBjNugcf8Qsd6CmHnVwadoCvxt312NmErIg9FnZbE
AM5S6NXz1f6x14ywC1yfNtZYnnL8zAXa734lgBahtTXrnJF+HjVMM5XtkNUrWE+9
0063yAuigcGCtAK+2FnayU7I0YvKZ3q7csCQn1iMaiD5qsarxGZSGp+WfqrYelRE
ZA9L7uuVTOnoeu2wZI+O/ZdwhOuWiJR9Gt+M9JZtTcA6G3Bm30sTsO23CeMNfWOv
7ll8MVXU843+F2OQq9lyUWD3o2P9xMpgYQpHoXBCB4mIRr/k1JvaYU/nzyi/0NTj
CtF6cb+WiliX4hTPnIdGgXWr5blKnhyKALYqzWWsmjKgfdc6oZn0yjO7My6KEBnm
QVBXVLYIY5FeD4VLwG54kOYeLn4AcsTscGUD6gJwOF8h4vjC4KQOEitIQq3DLy3b
/hlj2u8Vt487v7MwKMFg18bo3bKxnI39eniIVedhJ7HmXTnLo3LWH/QrP4jx7666
JStWZ5vC+sQIHl2LgqQ3YNj6y7WM17EtUtZzZUs8bHz5GgitSdRpLGcvrxH46kIB
KsU++SZeFUAqlXui3+7CmpUhQ88nQW3bSa0GHtfYEiGf8zyYWqa31s+YpT4Uym2W
2ZV1vCILGPiJ7/Hz/SWDZ3U6vtXcHRSlUJTMPENqcFvn4Co1zaX2/TVnTX4OLQJ3
LvgskkuwcWDq6WWkvCl0Bkkb81QZ8i31g9tVniNJ4ZQFjOA1AcB99ihOCtEH+eu7
Itzf/YHSAsliRgfKL9FnkO+3np8JAe8xZh8IGwJ2MwzPtl10q/BL8ZlVogplqHhI
KdGiyNKJ+09J7LqXUjz5S6qFQ48HrspC5LalONoXPjRzR40uDfu0i59FZ7JkraQW
6Ad7mQlbQ/1PklFuKLeyHwfamFSAt0FzvLVL8srTjEXlvs4R1pS+dGhGALsTzKiU
Ral+v+vmm4kFTVCnbWU0pNHDCYW8gUHyKejND8qzK7sXB5uKY/I1a7HG+McEYGaY
clpkEMWaBuPmqJFCTsZmWcWJh/1E1GVSueh8BZeeBfk1m+b1P8wSgrdq+59lxLhI
h26rboekZEtJ6KD2k7uDxY9UWrvYyldT/nXhbPIq1wGv/cTj5NxN0HOGvICfYwaP
nK4M+TpQA3/nYPU/y5fECuI/zqert1orOFc3aOzonHyR0knkM7VQQ9ux7tWGnfmD
v45NOnsNHiqQJ2NnGJ4W0GA9avWSZ7cQsuAvJTA/qhHrsX1tUnRg4fAclNR4EIDi
S8CpReS2t2Aabmw9d01jut4i9TFr4qPwzbDGpGsLgyPw3JnBDYlyAQyzDS9YE/tA
WxRIVOSmIBAnxfhAOWzPIRiAN95gb73AjEAryLBSCAxUkX2nLsHDuW0OSTFFGRfP
kIPszAlDtoSrvC9Z0c+a7q+sejdKuoKtHFt1jN8PPuxBlaOEqdBmOUQpsqE3KGiC
TauGGglqGSIG6hnplCqKJfMK4XzAAe7uuTXzR1leEJQQtStxPXTODFR9wtVKMM6U
QtWyKW+XcNqaphVtQXUJwyp/RozuX+LxAvJ5GSLKOF4ynF/yjgZCZfWgqOlik6Vq
ps6Lpp1bJZk7pGMgMsVvdxWTTaG1qFJOXqXeMBMAcPod1784m6R0kR4cTO2qpSu3
l8P/loQ7+FRB1QvTewX3d8KWIYss5udvc/vOp4V/Q9jK5ABBOtkLJtnyszhh2MsQ
RXngpqUMfDBMlDcx0viYgFjc0l005qN++iNHRXUVjr7OuCAcBFOlnW6TWyzm5e2N
WsdeFtGCGRyc4cNMVONIgIDdE9QTKbdfg+kFs37p/APzsGnZwckG1wSBKYCu4TW/
0TRoROwTnBEaAh2cyIHl/kkMho3eILKaVIEanohZ6vLCY/P5QOrS2v+sWAg/YMN9
iL81ydUPz+4v9KNbgqtdmbBZMp9j3Iw3/qWYRGXa+o3JVM8iiq/MMw7X47HxvEJC
ag6R18xWuOgbsQiHJq36E+jvzfgVCIEgQ9mmzf4fledsEKGTOnyQOKAdw2zXVf8Q
7LjRSPkEOacp1ep75UMtpxnLfJcatZxPThBWb2KGFsWJwd+VvxERRl5M7qToGR25
GOFMlsF6XRktYTx+4DfBWaJZt/v8KJrSLXS4GRmHBISm7b5YHKwBn5kE6zmF0DSg
Y1cwI1K9F5VO2Rbw/S9s9jw4O+asuCQzoZiaEvHRWTR0XdyXIX5N5mhQjoqIJ2Z9
up2Ta3vg0NFKWLGbN8SS5Pdzz7UXLwuTWd0cwuQ+8YUR8KcQtonahN1d8Y2MYc30
WPWNEciJcnw4YM78JHWtaQAeskEmXyA3CEMx+g2l/4YuinGr+moCATsrDmU/UBuY
pJz5AcgYTLW+a6ejK4Luux8QWW9t+CR0ZtotL9PhZ6SOTPQknmCBDm1MxMs0G9V8
sCB0msTh0pjQy2VQ+hRG0yzEM+Cf5J1aL40NWg3+Oz+6VHgxyywXxgDwnwbWCHIz
cHjGgKxS2hxRZ6lzx8OpcWltoKqK75qhexsLxYBGKvt8Tp9rwVA1GwKRHGDfFRjG
rnDt7diDbGmSxM9FGKRkT6cOcQavEz1azRK9IOdfIcd5EV3KSkp7Fu5cmmZcR9Av
7YBUmPXr0+5tx8gUjhxJMl6B5+0nQBYe/ZrPhKCygyH4dX5pZzOT18pk/4G+P6Ps
H7B/FGSMPoutcKOF5wr0fEsTg738IL2lCuHfjzw50wWT6BvRV0JyiGxmb0B47pF6
j8PkxItj7bF4qJBVSKUc/PPYaSSHNREobGXZ5bJo7a+W/uD7BkCVc037ioZlJRso
C8NqfWj1OgUpw2a8t8arGffG22Gf5TvFdmLN9o1MUXW20DDNeDUcseLpUYDpWA8C
ZXUl8s4OD7exWYFTxnvEEfd7ozCE5CGZ7MdZMjoJmMqz/UHGWUJNxE69oy+GREuc
JANSd3RKiSnV7uRD66xjz75/RNg6c8OLWdmnqU4xGCZiGYvgdSkaKgov2I7SSmTA
p1TXAT4KFL2kXO2VwD8M+eTdaomxtin2TQN7ZMVDLV6Jz9ie4RahmpdJuENUQdxc
hF0bgsvkzCVd7Ya3wvr05RJNI46+k+dTCpcx2i7ZXMIDor6rVyAjZsvQKIMMl9qS
ATy/CXqNsVUJ4wPoz/xyaIkbF4rVfvYOLo804gGiEnGszkb4XGeHn66+sT1oehBX
3aTakLHTU1Gny7i7I4J9TXGs5tOI2KezDrEjj91ASXb+fIQrCT1qfwkXt+aVcw9g
NITuRW8gCI+daNVhMf8j1pzj4GG8e0VQC4508tFfFiuDUoehpyehVUQ6on4ma29w
0Oh17WnjWwbA2V1NaFKJlz/rgZ56fUTisHbEHwkIb5cKj5vnDq2lepDdpXosUTdF
OiKL5IOcgyJxIAskT2BodOvPEdJeDvCcq5+9n2+pQafah5blbPvoZsTuWwQEx0bz
ZROuC9Stoobw6e6gjvJW/9S1RCGGUrlyLHEf8NxYhqf4/hw68hyYtHtFQIdR1GGW
DiMFCg5yGdF7ZTabbLVY/ZLwAolx0Fp1heSC4mEjwWKdEO+LNWBg3P4td2tRqqsj
Lc2fQ8wzpDTIK35eNRfZrD28OorCVfjTnJAd+ke3d+lqZib0Cht4XMR7Aw02Hqa7
0uci1xT7hSNtpQqgC3sT0Cf/Zfoh9mOD9qjBUX0bG0sjVPOBSgFTTCaqR1CbwVJL
AZKx9JOtDfTLbk1HLNRxxxg+pOs/yGXCUShNE5J71J4AdNSDB9usp415bKEmvbG0
obX3LScns27z8fGaWXwtnrG9G05i+y3kgMIlY/fswdF/lE5O4FqKvYJbwJmX16aI
k/yvav+wxd71e37B3wyZXtNZ1mCNuWBh+KArBJJmC8X5nFSJ4qF2kiro/0g/sBPg
8N4iqtvdm1cYeveh3p7uXsAJDnEljsUkMlrqq5q6EQo41ZAY9/UZvP1XFZghRKr4
6QtKpKATHZGNHpnG28GWo1jknQkiIYMUyaYrfeILVhOaJL+Rt9Ua8zOl0Di+ka7M
NTBG//yOXkTBniHlKsO4WCYhFnFTgkPF0MkPaldYUNDutbm0N7XYGXzQHD8XHn8a
roPPvf+YVOr2B03XBuc2QmNVCcAR9rpqo9H2oCSBb5BrQyXM6cIWdjQPB/9TYsdi
7HYbIXvtCpQI34obqChSugbqBxvMW5toJJpk7xiugdS57LLllo2dJZGseoNyq9xY
52TeqxJUY/tASY0OLzMNSJpVs5QSK9S6tC/wPQ3Lb9DatoOeJKAt+gpAWzBqSah/
ykhsWklvGpWcN/ti2ukk/OMfZlRI8M43zotP+q/So/FfGoAXhxqZEv+s52jWFrDn
ogJ3Wbh7pP1rfknXXUq/asbXS/9WX34/iuUUfczD7+NZj9ulzqLiVMQEzXp9UqH6
i6eT1nuAE69rf3C40QRcIECIuENtpP2fn58UdVc2SWWUR0d4Ss4JFQ3GFpPduJHO
hQ0aVwznlZq5s4ZB0JERQ1WELZnMcXiVzL85losgUvK9w179YCfwiqsRAlRaGp9Y
4fSEkw0hDevNUgGldAy0Ft790tHLOrqG/2MDPZ6y4cV4BU5oGB4JUUaYsFs7TIxb
VTKTjEoupAmaDG4CsIkjCoz9mrRNcG6l/24S5GkY9aYVOa9W+z9f7FGNCAYnegXr
sw8sm72F2E5zq7xpLfuMjrVajqEl47EAJO3BGj2ulyPmeTyTqx2J45YKX5x+3MG6
vt4wF2+URi6SkB4+7ggPlfsksqseTZ+aR5mK+DQu+J1dZdEIdcn4Up6Sbx/ImTBb
cUNafrAZixhOdAfHYkTUufO2XXxL5qqGBFcQEMPQ0YTiFU5ILvxTpeYU3d5g8CyU
ygZwTmlr+RxjMhio+GGA+qo/UvWcsojLKjQzKzpbg4N6PQt5LuDMg9xYaB1lJcq+
WhAZBmB3F+lT6k7PZchDcicC1W/PLLGL+AjpntrdB/3x8nZptwORRe2LE/CrUBLM
ey+DiLQPPBMTqAOTYEQiSkLHyptOzCpM4j/bPTIadfb59eSWaD1WncXNN64Kxxrz
/K8gUv1YdlxO7P+bPz7AUKvxbiAGQCOdnFvwkbV9dkzQ0IF3XdEKgs0LPpmWpN3r
R3y3OzQvSzG7MyqWTRFGwQ1m0TNF9SJpsc9VaYtehsWqu8T+s6rGa38rd9/Qt6X/
C5GWc6pr0I57Z94S2QNg8SRm+AGLuBsILdqe//kKSs7IAkPnG9SFIeJPzdPjt8m9
C1Dmv0UFOz2841IQjBemMsUnelF5l9jnuF3D8nBFCRT06ME/L/7II0bWj1AuX0Vg
JAV4lNEiHsBbkNwIgQxzfysm+BAP8oOs8sPkmqDCl/BERTTGuxWkmyeDwe4x9fSF
H/bmjpxolcYI5nn9u4xahXUiYPkqVTc2bbx69ZNi1RXp3RmKoojeijI3mIwzWvxS
LuA2p849WrF/ccYKust5fcRcwQfl5kxLMYlBg4SocGp0boIKJXdC0oaN7eKi0b2K
ACOh3uP+VAzTaheMIKRRITNINII/N+LEw/66C9dRUayL8FClN6jBbscSlO4mM7b7
w6ZJEsRnc+FfPlMgjxBYuNWKV42IzZTsZRXQE/kY4KxIYt4zej2iC0X681sTe9vl
wi6YPBZpFlubu6nsrTIa072R4Amy8V5xbtLE/GT23/WpexJiUPjqicY9Fr1Ds7Hs
SXwJ7yxN8QSOZYTszeOb+OSGRwDzfyfpQRuLLML0pVkw9vwk3aBjg9bbpG5VEXzT
GG9/vsupp0HIzRIm0wBnnHVV1D0E9p+9xt1xmTRw8eUiYcilVBeo8Ni0zF8iDwzW
R8Q+ZMUKjQO/ll6d51ZRc1jCjakoQNRqdZl/aJC3iMNKoTslzXB9HNn3WDnVI3Ro
iP3qrRjIJtQlkXT4gt0lcgaGC7ogsD+bD5V7v0PPkVme/cwNyevUF6xGS/m/fm64
ZHFRI8FOhvL6bJkBzQoJ8ULIKsyfWgiV6HQcP3/GLAVr6g09/zzRxITouUGV2nIn
UO/j0bWRfgO2hFKr/0jMB2l3g9zzQUuSeytRfaNctTPMWQmD8smwP0lAR5fVe4i0
eQSpn0iTue7zbe951Lt3ucrq4iQJ3h0kKlzwJgWb5gw999Ax1ffnoMGcyP9oO0+9
7iicIU10XRBNDCNdknsNOC+Po4pi9CXzh0FGEEIrQfm/GfWWF23R0zpKdD6jY3SI
ixBHoT1jbYrfmXseypyRp1mGDmuY/9mPn1Zja/vw5fu6vMsqIY5UEwJzlm4d65+J
Ayfig3m1offziP4pCHtgNVe2fGDQLDVUvugqDQwza28WWs+CBo2my2uiXo7XMSHP
abI5ZqIJmmIvPmZgY+48y5o4VrdU+6xhoSlNv2+f7rV/+/6qPHl+SHld0+GOdC9c
r/XeLuFCL/9m3AJ+SouxX2QctEAESXlBaFuJX++Nb/mnEq73Dq7vS4+SS/K69aFF
r7KWtYEu/Dvxy+LupsPvJ/6eWcQcVPXnkWBlN/EXQFIdOIIGdZBckjWR5JMDTt6l
1at6FNZanY7BdQMr3vnsgzWFODcSOab5SyTvpz8ZCweXWwqsJGquBKGTH+6T+ALw
tRggnyR1zMYXdJKtls9/Aym98agatRhLeSg6Gor/hBCoh5+wELGoaLpGJhRuT3le
YQMJvdzs/bF91qfjtznxbXiaf3Z28fPJXdCAc5AmxNEOhqg76YdAiiIL0vOS03e2
sAcR9HtCE4iJ72sGGGiEhIT7R6t5vhE7T5K4NOSu8G2cQeQ4bf5Pwxgz4G6T0QwV
S893nkuwMeQ2WEnson2UrVIOFt9Pz+uG6lyn8a+u8jauHzug2jZ8ks/Ehx9UQkPF
cUPHA1ntdhuBFwI6IU/ywzfyO+eSRpBLl4ake55iRyzAcD5h2Qmhcc0jMASULO3v
lR+lO32sMGaV0kOVhizKSICOi/FE0mKmQHa0Rivkebq5caTlwWC4MTlytRz9x+Bl
FgzJMpZtCQIq+FE8vfHtreZfFJpdtQ3NZ0MiYgXTjjerorzBmeZijLd28+P6Ghwl
QMGXQlqFrBulFcFEWBMRccParNn+LpfawYY8Mxtl+LaIYoOPMcZhP6GomX2Cn/gd
g5upysbObOD6stbcHrYe0GapeNq9hHZkdJlZTDQzewz8CqDFHN5rCNvxuhS1Cmvx
GTHQgPtOOG4rxbqrAF5bLimyCWvWHM0G1eebRUSqZtGEdQzxwYAl0jso5JCZN0IE
yJJsZhU78Evefl8pn+YgW1KO70RUqp5ZUA/6OY6epspG8ROvLlNTf8710u2xpdoy
cKmlevUO25GAKQ6YCiBBWpSSZ/UeChTO5P+sxjI4kAWX/e7u5pqmqUxgQCWirJRy
qFXFr7SAAp9h8rGHW2820ErvQEXrBT84vFx6anEwkvaQbSj73Nke+qY8MZGMtv6h
hGN9Ohr8EoI4bAzz5AzLdD77ZRKmcnKhhCqxSir1OHeL+LBc5NRSzBoK7l/GK+Ie
dQl4Z+nSFkaHEUjlc/1FyiQH2jT70Rnb0PmJL2f8u+shbaAMfo7dy5bgTA7OescC
iSCYjPUgfXSUo+k8bHGQ/1jL0jajHMHpKh18g8IVqbT1i3PBjCX7z+8Y0gKlQNLG
91hxExCpQy+mNj281w+WKNw3vSU+ZN4X5aRJuiKxn+GqRj/a8JyPx8FB6V/80q2v
KOodkZKqKFo48adQB11OQjyOMYYvDP+aymY1RKrj+QfD6fHPcEPXrbLk4Jqy+iwG
21MyKu2UKv2AJVjgrR31eunb84ZhJUhRkzn0njn3AnqWV/VL/qkUtbPdHVzuvYjF
5xJArooULv6/XHaB9v5ihX9vxreUSXQjyVKPGQuMBaW28OOqg/6Ql13bty41FYAN
gDzdGpPdMTe1Sdm5Ul5xtu3Hv97o12Df18ipHxDxAjbCQ0b9e2t4CA1oQCUodADQ
QDEBanoNQw3o5u0P7HdG3Ig9/W7t4oH4bun1kji2dTXvUDvYFypO3yD0thBP6F3a
DQGmwq/rcEmBLBA5tFl42XoFRNrhp9DmL3CWY+T1YO65HI265UEEg/W/ExhLeN9R
+gbq6ogxLQxKCxj68qUmkjCFq9LbZvpgOVqwpfA0xXC3QJeXuO64LleUQWM9LcOI
0cVY4WJI+VbjoY4T5LfxYezZn62ssF7HAoEP3zZ2QbGzqi1V0yufNad65X9HHKBs
BwKRT2R+Ldwn/LizCFR4o7WLmLpre3U7TZzOWyUdY5sKpfvSs0G+10WwDvgi+pXh
2jdcJTM3DcG4v+MmxnCGQzB2YqFObx/+rpenuYNt5ctDtLStClEB6JBGqq0HuzvY
biacV1k7Yi0a0ymtArt+xnQKO+MtoBqeGdMNe5kOferpatJnb9vpcTonEQDukeY6
bsxW2HL/+i2GlEFniGBPmc4XqD0ixiHZBxe+gXhqggfEK57b/NMZ7hJdiPBFo34B
QJCTgjt6Go8RvYKxng4qIWHORCbI/NBqQb36bn8CpZuz4ZWi+G4CY2h53YjEa77x
PbwOIH95VmTBM4XdwyaLL0l/7Y6EW35LTh4q+kMktcmkO+K4wsWA/9aM+3/Tt9Zi
GhrmK6Kze5nEYEfJPWjKuA6hmIruiXgYYd+D2oJ7cCiMZXMRk6NA7aeaNGo2tauW
MwPn9KoBAosiXnmGmqnUY5zd9D075aRTj3Jx2EdOc+wPewPsYi5LFVscuWX5FB8T
Bas9y1rVR6H5LIIjpmfSFoWcE5ynefvkjUMaHhnWtedNZDZB48OGtqbGYeBinsHt
71KwFp+Xetv4ugcEW+kFIExGIsMkri453Pz5voHBQtZgz1/nw6w9ePOXriGQpnBw
QoDB+LI5tqwP4T5V1ytDIv3pPUUI/4pgwqL9SVgEkJKWJrOe+9C/QRf53sQUcXuK
T2zjo+SiCumFRWbYctdb3tX1LA2C1eZkCryb1H7Nx2fOPXqZTvkHKBglvZ19GDHH
Tj/b7X1CR7lfiaTHt60F7Y2GbgSBnUVM/Qc5rJqpdSlnkJmTY0IhWSp7nUiyTyps
UiDEr6O9wS09xpvU4OJ4wcT0hS15cmVCnIjuzFaXSgSMHhrxtF0ZShfD5qfJIUmV
l8ixr+KvhICBkyUobRV++rpb9KBtD0hSljv6DowTY+iwiIXQJIDSFaijtHhCkMUQ
IEQnSFTsIyvoy2oXaGfT8AwTb7bGbDwdi3ZtFagl//954cGfjMhQpdafpYnfOeCw
VYc6iK0H+Dz6cKx4/ihu8RdCODU4VCDTtQWgjb71zWIi5YRIRAgINsEbc9UPIdaM
GUVgeB4nAvZ3/2Tb3cq9dEzvzdd0pR0teR1XTRK7m09zCx4bM1+R3SMydn8nwGhT
qXGBKUEywNTTIXO5aQTTEqHSs+xWMuZxNQG+DsveAU/P2rLcLPM1rr+/cJpWbfLZ
Fg5g/rwQozSLZ/XQNGN6UT1PMte2ED92NcopM2oeSDzYA8QeR0LJc6vdByVLIg7k
rGxgSMQGfgpOVQRZk0Gq4/1gklPKospT1kkrPGpC0sHcBbRFJZHqlR3gubifT2cy
nPyt0DGEpNavtDQwHYsuIVdN7eiXGJ6sl8jQKPmnqnQpeeBR71GQrf24AAdEDJZQ
qn3QdN69IuZDXT5nAjHJQ37CnFAubijtxX4ZvJU07uYbJ0eRr6Ch7rLfqWRaZSL/
ejINYVh5N8WO+iGOU09U5CBwZsWmQuPbpljqb3G5pByGcy4SJnZPv/7V/nUQc59D
3aHRT1yBAs4EbpyyhFLmaq3KB8hSmZvLSaEd+gUVMo4VuS2O/XUX1cAg+41Zu3S6
wIdLA+MFvZakM1rtuvyyLD9QHw0rJXKM+7xVikXMxb5sDyjSMFSLJOHrIYsN+0v+
+2z8BZfxaWJTBPbjmRYgJDf/SZiX4dzisqFtCWvSs1k8auUdHmo4m3TMfiuX7JbJ
gX3T+EWPmfaTB2W3ZMI2gNBXab6cAvJbna3cCkKFM2zQD84QOJoeAbZ1WvKAuuTK
JPPyNPA8g9R+eCii/0rsLHV1L1saP4OtjnB2Wlu6Dtv7vgezpAagHD/rGU3Hg7yi
sIGbrtYSHT2mDo+BeftOFtEQ8u8qFDNt1rYNFpdv0pp0T1AFyfn7apiamP8OcICr
rCwFJ3TzR6KHbpUdij/g6BxGpT+5PeSBJlh/OchqN5q40T8EuWSGSRVKyixg7xyq
QXwhUs4RFwuzhs422oCb1MXWk9b5QK39myS8x8wEzx5Dmp3LCbELAAExalaT5oPY
zPLKRnZgnMli5Uzy3TJqk+l1vbfTVNUTsqXOUGpIi3xTNj55pdg1TCDwZLfMCYcm
NYjqoYuJqKw9O6Oy+x9ZcztIMDqaUpziAkb1OLrHAe+co/AsmXvK9oDZLnxRISqQ
MqVjNPY5wkz+OU8Q46FZXnq/+AzJhiGc4OL7/7P4Pz+Sp29OgtvMWl98249kdCIw
TWo4yTfFHZ/Q+HEsaLFBzUvg05kLvbZE0dTRERScPD+ww2pstrGe3B1oH3rENiTh
3+2l7e2JDGfDoKzUTvOPsX0b2F3weof82+YpicRDSOK5V8xgILhpRURBsJXmeI+Y
AJxT3IYE4LWwBSpuf7S8wMvcOlorLQfoWUOxsvA/J4dONGdYu+A8hPW7rAOsQMY0
t/uDJOIPtFBNg8nutiGEevtxoVb6zTsucvINzYQC3jhJQMDzslYFrCqYDbr/zH2W
F0IL7Wzp+wyA8vjz6zYTPEpIcjavoh5WvIV6KVWeymcHPJ9o3+ohYqBRe2ST4Vp2
n1rrThS9s87LcmPE0yGfkiZY2racnHCmXw+1xe7q3rtTnhNhxiR4vCdX+7rlTXsi
elkst1tVvTW3012a15WkWkZIDVqxG7rGZ79TzES+fc9M1y8rGz7zcXJJnkRUmuMZ
kcDCqE+WY4V1FWjPVnawu7gfLCKwnGmk6rwBFss38oGHB9PgvcZNGDn//EuQDyGi
wkIH4T7Fd/wFPTY9N1X8OuAXda9Ngjs7wqV7Goptk4usTF5vgSHM/axTX0WCt6Oj
ZDHD73GUGgUhA/TzdddnZowMZCLxDA25Qqd4uiKH9U6S9bc2eM56LgNieFRmXZLJ
DCyt/cydVSGtprJn6W2sqOfWZlKx5eLzPenBFzw7vswt1aT1UbrS2TEG/0kJuJG7
SQ3OXdInuvh/HY45dWeOYkflphOHox9e3W3OGlWiZ8MX/5V5v7huRHfgdIMbNcCp
+MqqNp2Ykt7CX7ZzPhKQyzFeB5121I733b9zvQCwM3DmQZydPJRES21DDiSnZK0E
2NC3BEqfxiCe4Kg21v/vHC7iRs/CARMU0dUrOZkxL8FqF6IOUuJmbkSJgmCnVNMs
t/RNnwdO2npOk1BG0QmASjxz17ayGb/xtoFP44ieCJluxK55RdHT2FQozQ09Ujv5
vI3qVOj+RU+5AKPPnmABcrlDVzj3wU3eO1tgc4Nd2ESKDf2iSjacqiSRrA9+Xdca
/aujwIHyWxYXcJBO4HT2WjbhhE6VLk2sXfHSA99XDKsclgfkAXdkcM77YsgB9Lcj
b7CoZkDa4CG+Mb4JDvUeUvBVrwingsN0msD74uhQuOh3MIaRIQ7eg8aZg7BGOAbB
R9Q482jlILPOge775YtfJ3vHJdAWJqFJFD9UuGBYXHio9wTPLKvP/m1FSEBKRG+Z
5U41Z9RUUzA0jAPYWbIyMf1i16fAeCQmrOSITLt81a9/ftzXX5ojFcdkLgkI2Czz
o2yUvjDXI5oR5bCRGODUQIJ0XX/nQt0v3IR3HIAfFyjdBcWDR4C2vtj8YCR6/Elp
4djKC1L1Cc271MSIuGlB1KVxPyNYT/XQEM2BoNgHavGgRCjQB+h/DlEefR+l26tx
29efocioKimHiO5FqB6kCfunyTjuPAkQ7gbO6y44DrgLdbHa3TtBZWTuMALnvQdp
jteU8bbCCLfG54sCpMlDo6J21zyi0rN93JDCM42pRmrByh3YBrzmYg8gPxvoKzJR
Xva1Hs7XPG6rBjV46toTrcC3PeriPbfIOyMCyiihdBJZjhdkMnTY+CzQqXAMwlLF
7Nqoawi8T6hwqL4KFQRoYXxg+AU2htT6K0TpR6d2ZWeOJHZ9Qry05y/s/ITp+S3I
T3ZyYckPWyj/Vx0XalpBrPwbZtKiGz9ZWOx/m1LA7pfPSY6lB9KPYUCYAyqFsEn7
BOCHphQoNPH6NegsY1tAMeuvqKp0zBmotn9gtkou0O80XuG9m5sPq0QaoHoK+yPM
kywpnkb6jsNBzrLXoFHotR6RO8quadyI7hvpFIgXmn60hYAg0HHfjO0AG6YG3T6Z
eighEsN2MuBoFqJ9WEFchaSlIp+fmqLwgZaqYKAx0WAoIPzOeqjt7yqlYWZiBEBQ
Em+hGkG8Bmf3flg9h/hX4YInf9iOz3745koGRmig+Be0/VBbDyuiO6tolnuLsQiV
yBaUdTNY9as9Dp3YVZ7f4RUa+PraIR12xsbKVFveYoWXcAMlO9CWNeB24XWGnMtW
AZWDkhoQ6rbHdPdHzL6U2vxIl8I7cWGhRZUnLcAh9Ltz6Du1jYyazmTeXo9mE/1J
ngKrV/rmeL1v9hQUpBriDVkrYZibqro/MWjXOnFI7zMjge0yCDSpzY26BVckb3HN
nFW2jnU3DmTDzX8YZCorAJi7KdMU92V8sEtIPpUnhkh6q4d590kIYHBf1MvzPE2+
08P7wG6hd9MV1lT+I4Nqd8TKo7FtoP+R9E9goYkF9JCP7ItUK0RJd5TnW2JWJr/W
dtbdt+okCGDui9ND5dMLixMlX3H2KLR97vEAvnoqHrfhQZTb4Bj7wIUVq+BYDOhl
qLhna7FdrRFCqiVZHhzfFvERFi3HPBCIztU88Y2jfL/vZuF2bXU5rSOjU8Ht8MsL
FFemWzSngAO/5czv/xic8tnqi82QJZAuaE9hJgutuB0DsKmiCRE+rnZmaXMlRFXN
Xp6XzAw32luo8WHgHhvIZfifYkCS40Dx8YST+usBq/uwMru8q+xyKxhqm/4a34YA
mo4RMMQ7DwDXLqAAtu3JdZBeBSYJqTwQpCGatqjsh5RPLPHN/d9uHjnByduF9LR1
ENAE/EfzfMRA44QN2teqn/DHdr6ODCghCJZ7bic1AYVFRzMVV68vRfDxelx+tIV8
1GNmgVLC+lqPY40Ii0DFeD3ZJ7dS/gOe1WrdF0hVrbmW9TgLJ6zSg13GUa5P4v6R
uG6FB1CTWfR8q07l5iQnIYbj4YOldQZ8ondcts/iitXXyEUCONXyOYbrE3S+Luuj
un2c245l2qybhclpvBuCi9tOj0rzFnAs1/sYXEul27IMDtgEmKURwu0wszlkzdyZ
JrxwLFIwMgM1tyF0sOKbZKLSDcpbKiZiSy/4CnD4eYvkSXWy07GGg7HXxzM2RDkn
TDS5E98Ajy+mWKP4ORT6qRmFrsb4M9maNFqXx7lCHe6bGcRVm7/eNbLNt1ZQ3Qax
/FSiCKmzlIc0L82oordFDC7pwGqMhhxcnUVyQrLmS5LSd6uVHXjx1SEVMNvx3BlR
5TC+L1uEDLpJjIraQ+IODo4J7QV08t1Ihg+NDkNm9v/w+5M1OgFCx4xzVd9IfSqs
OK7pCR23iYf5pTbFNP2CQMFSe6TKF3RGO4xmyCNCyIuECVkMV7O/lMdG36gaDxyp
uXNIuy4oigDtH179+sCHpd4/dEv5owjiEhRjy0dTCZWvMG4O4Pb8i3amJapl2uBs
TyCTRuJQi19Mbk5TzVvaEc88ihmrBwYA8gdmcltCQEE+pJOOVNkuPfLX3GzKD/Do
bEp6z863M2Bmn7gQ43nibp4ZYdDsNZESibgrG9B0JkU6U9WQDp7agn4hqYnuHCan
31gUNHYlf9g5FVx+3WGGdgk/htUbNTr9SWvahTJP2KU5RF4/Gx7M8D66KF8N++bY
0WHeH3Sv/pDs+m+PeP3MQXem7JCRn3zhPF4baWPFzKiL+8HiUuxakFzuV8DAmhhf
xFVSjxwGmc+ka9QmMFgIADvxnKPsox19e8QlLodbNdyWzElpUgq/Ll/ligLh9025
X3dWfFaABHGXDnbSrq5IRwYPIXR71Y0XynP8hRkfx6p1Md+klTlN2miBNFzpsBtD
HmPmrlfDLnwGYBYOwmBxaI91Xr7kNkwYfb+smdu5vUbxtojCJxZeEQmlbtEgd8cw
iS7c+rqJK9Xran4kpNdllsNaZqddkUWVYqxD5Cc9wl+lCK28t1Jd6awjKOU6jsSH
P4/uXRjnZRgWnHOqxJqFC916GAVLs+uAKJzNyseLX1YiWVpLS5hcOjWdXxVVAR67
4rCxVGPbrKlWM7MRpRUgmRy9kW6DsD6rndy1GxvcxeEiXrbzwxI2k3ue3l9z45id
ufwX3aKylPuuSEhJfIf8Tj1KyigwAD2Fp714rj/3I5vUsqipsA94K8DcKTletQfC
9/t2NbkHu2czr2fQvRRUmEMIK+2XkPWV4q9mkr11IqxFlBfBcDWZ8v9UdDPNxiUW
lsFioyX0HkQM6ACLvszvFFVmJg2lANRqCRNeRdnpGNB4j+cxADlTBYo7qAot0h6F
YedBS/jrgl8gY7O9Nfk87TJa/wUsA9k1syFRQsmjnxSWCUduFDzPBbtnEOVxb5wO
KuFuEi2zryUiTcnEWS+zpQiWZaUssQRSZCmunQ75TfhN5hPSPhHsE4wFgL+lVg3R
IukthpHElutVrRKduLyxbQfFj6us8YqgJbqC7ZLp5q1J1ZfA5pasSkOJGwArpaXK
/VXAWO69aGfJgM3Y33bJqPYcakHWbF3PVwece7qj907iieQMKoF66no9aZ5p2oo9
ubto4iW5TO1Yjdo64O/eaWXcGQ+lDmL29kLF86tnnvetvpSDbG9s9NTu+AtS2FKD
fdkvJgLw/ZnzSYnNdkeTUum2nxZ41IP4f6dSfQdSCLfoGzDYyBPkTk0pWRKgSvTj
wvUt2fsF/btwoM3y8sjeH+q5YQ9XhNA9gxWPdsFQ3Cc5lMEXjf4Sc3GzSwT2SaaP
Lc6ugxUCLJVCfyNkZg8Knpbkkb39Hsv/yGHyLlkM5L4s304FbBxWXvo0OKb0fy7q
CKlnJbOVQwCRf4cEJrF/yyAuK23L8oKU3r9A0EsgRd1vQCI9O0PAkU12+mFoYhGM
khNZQNPECB+35rPGjDybOhN8en8oWv0h+++LpA52i/RSvV/5enGrwPjMDeVFrBss
n9xupaMVsHxxDJV8msvuEr+Rkff+KH4EiYT7habRwhqFnK4DNT8hJoNb3oBMn7Ui
HYP9m6dHWdtf29bgxuR+lr4o2RGatKCxXVJNIpl/Fc6brE2gisbeJIsN7twB4LaK
lT8js7CzWy2J15xZiW+mGo6rBsU6Q+j/l6FC01UyOFg8c7j6bZeGXJZZHzyy7lN/
xQMQTB7wbokddgh48QcBS59hqBlHUkKZWS7+TGXqzFrPOToHWjB9bLnh2c2olS54
0LQADtpVUl18LA6BOVjhjLFaziuE0oemrZ1+aQGcBiFARhXUYjH7AagcLAoeRmwd
r36mdz1E3DDgXb95YVdrrYL56hkaoUisdi24P7EapJZDAdkp4Iuw2o7JQWWHnnAG
13zczJ4jE/GQoDWqjh4llAVNuzwT9zndDLWblaGkb1K0q8uf9uuoEqJFjrOBeEcb
/lHb0tO6WH6KIm5aIYuLnM/AOhNTcvezVpz9jwqhjZOD864+IMStnucA/F5+NjU7
VN5wrwS5MfOTwX7bJ+exmPuSg50LY+NcgkaePRVKgdHY7CiYD1nKk+tdqBbD9Rs+
BHjEa5TO/tJ4P+oznuGKliQoMTlHCshzLLj1eldSB5SkPblF3sBc4MEM0c1ISYda
iht9/TnXuPjaslI7mv2vC5vNPMLqe0UjSr95xTdnG0iJFvIbJ9/21JB3FLqvmQHH
Spjuz3RwIwdAjIb+eH1JxzVrd2cl8dZWYCfhiXQEHk8tjezL1RcqymGWMvCuTN48
aWLSR75K4ycG7heD2hXCySQRR0vjNW4GVPPNGsHECQhXOCepv7QNH1KyR+76D60J
dQzH+jc/SedjEYprxCHBZBI1Gfy2nS9zbL3P03htJJ8BPD7tqiIwhUFJPzpAwTqQ
AEE3Z3i0r2CTmx19nE4YApUZS7cJ3IxIIM1gAxHvsdMFnOvrpEAWltRM1RoYQM3o
yxLtsZf5RgNSPLoI6dloOvvMdQp0HcG4cnM//H9YhUDOwdfhvAZHVseHSN0e2sFY
Fc8QS07iN/EzpYUZCHTaS0iZMigCAVaDOWXZ6cn59oQUl/yI2gxB0+16SnXL41Nw
n6GOdGu3S2n5x4lHNt7DmM1ZYBsoubfulxgg91U8pA8kjf6vn9eb9Ts76PqhfxEk
sYj8ssfoAPhumH/Z7UUXEadQLQ93RnVFrK9HbVYWVgExd5TxUSIaObFcxqOLAIW3
lyfVScxPZIdikWxRYzBOdp671O+wv7qiQEyPPk45fD4CLQMHslSl57ouQ5Ow/FeG
amNXWj0FeBR4ECbB0nkvf3cEDGeOpNkS5PTtCG17L10j7YGrWryYA5rJFiDNViMg
wo7/JpJvvhooZIeS2QCXhCFsWF8QuWWiw91DXY6l93k+lgGq1ZTaWbkguvQkwNXn
oZDOwVYWtRu3muPFR7jlB+78FphmhJ7BXdTaqGcwBRHjw1wYnrC60QoL+0iaU+yx
f0KnXDPPelZpHmz6QqG2CEwPp+CAnXFm/yUSd64j8Cyhi6oIJ/aVS39DLDcc/7qb
Qvw1qA13ypH2mT6j9mTH2RH5+qgjrYIn1uRpEtNS0sepeSxjYQKoHYUnRebsNTCw
7RxiQBBCyqzqWfy+eef8xcWKDcOePGJawhqYL2sQKucdBk/7RzK/fXyQJH0Ywdlv
G2Ovk0+rb/plFqArZMxWsW6g7g6baPcaqxz4iqiEHzU7GoNnYi/pIGOgWl/w46ku
ljaDZ3b1z7oA87PDIzehfwILayPhJho/ZI8YlKUqvacP/pmVQct7DQLpcXDC8taN
blpPLIJxvz3SJZ9CaLZrsrohs0phsCldYA4OduNcLEfuGatZt4eHXkYec2xslv4l
28c6f5ld7RbL4HN+QvFbli9saZWRi5lf7bYXpPlwThF/5dzCEyJ2tCLzt6dupFD3
c7XEe9MBy9lpU9FxR2GR+0xJHHEDS0BSrivN52381cYKEIbt/TrCkMpftfthvjii
SmFYLpvxTqFVKzaZ/XuGoPCUbHMf1K1mJqk1BNgLwzQObmqaGLyLqADr8H6TjT3t
9GPrC/87Hkqhc3J094jPFVDusE4tpWUNmFk1xU+zwXM9kHLRPOTo5nS1g5FYpMAX
k1kZ8UYoVPYb4Ir7GQS0nDuO/RjFMcA+R5/xYHw37xEYuZ7Fj+jSYI/EJ2dhpQeQ
0vEa/Dlcp0Vt0loXRQPzklljC7dXVay9O5om4DmlUcA6ssAIKzhCjayCGuTkW5Ku
Fhvtp53o4iKqGpMR5wx6O5WwbPOBoRwtpkdhhR+wL0GOz8f8D+6zANVISaFKtLZK
7INNbm/YJVDZu4DYIDsq96QAycRWprkgOSXcA2wI+ui2s1M1ZY6Rnz+JvO/f/P49
10FJfTUWQPqsNwe3DWpTVuPbcFcN06Vp3IAiugZ5e8ugbiMKJNgKjULojBUDWRWb
4wbYpLaMOneZyb3cymwkASOOJlkqBh5wHMDQsoiOgBF0jvKxxzwilipz7c2/LSbG
1KmkNThou45sPyepB0udevRRodPLUGsIMIbFIMhV/6z+JVmNxC53TpiDo5IQYHcQ
6XRxHPGzZym1LYNAjyAPsgZhOOOPcdG7QsFhSG9C4ShJuUF8AW50+J6R2SviBYyM
hfkBeF/NiMJxK+n4Wkb6xoXy6uAU96RbQu0xMyw1+zvB7KlBzJAXXmrDT/LvYGXN
ACD+GrY21Jsd5QHwiAz1LuIcsXHa4SFJJehXHs0PzVh3p5Qu8SFcSOns90wnfz+j
D6UxHIDwfIYE1fUsBClhfhy/LK20rJWuI76C+p36vN6KrFtIrDbysWgIPzWA580D
fQoTHpvtMTYFJ1vUlRLV1re4/XXj49FKmY5//GR+9j3BiIP1/O41BOnuWMmulsGC
hyCFZteSENUIQTTDg8mSl3YYBQ30Z+1thjj9IFABabREitDb4zWhtvlpGZ+lWcCv
uI1584w16213yYhm9sCdOvzsdILWBdpZrk5hby+uJPgzUBIAMotsICfwIschp9Wk
g8BU6RuDgbBjgqSHUtqlGg2TnrDUma+uwHUUtcN/USrR+PLuaHSO7lw+2S9Qp2aS
Ml8q4w6yeozcKLKh+O4Unkd3jcDZjPIHlWXdd81YOTlLk2L3txHcBD7Z/xsoPtD5
xpnX5a/ZZHrmvUnPykE9hXY8opVnFLn2o+8sv5p+Lusrech33v7ptp+joz8NvfI3
PpouKhVvaQaw3wWpzM+V6vEdVnt7sDhdHQrWu8CTnz8jBZMf+qC9kZtedL+dgRjn
4KusS0/mCeXscV84npWQ2gd1tQTAr1mJwWDe9a55e8HdPch34lwfTl9d1y3vITN/
qSQ53mfSwyZjCWYB6CLfHt4p/fgCcRGtuk8AjEvJCjUiuWEnLcB9MO/JcMyGLzn8
UsrSzmUk4IXoUsm4jv4BFy6rNWV9XUXIeOwjDAqAd7WXeFFVYIK/IAx4MZeMBKb2
gyW5Fx5Ooj6LsoHiXqN3MaQG8wPSaPn5XZf+X5nBSFfP0gj0GYILC2J7TOQmXuMT
LS0rOenm8wLgADLbD2ggjqMiDRgOkE3AiXBEhHeFjrHwPKYHY/8A1IQ7XfdmyLdN
RA0jeL3vpMwIoQrghkBPuFncAvBVOCVDHHt1qT+ifw0X4x0luOq1dz43A5LSU9ZJ
ftt5fdnjQxPjf6kBfWKGteXIi3++3vnA1jVRwFZzF0GtkDoJZnl8avyWSanGkwaW
OWyPwcp0t9GL+/08EJM3lZbnofNiVovVBnlDj80AOCK0SCaWL4s//KK3p1bGZ1MR
uEghVVrYzwMAuP+IqdcBByknsWFYk9CV6T/tIBN/kKziLLJ3rmHMYdq4yS5VBjKV
Miv5+YLZJmWZbfJYgZt9hwtFGVYxqFRBYyw4n1cEGdEF0YrEVLY4OhSK7jknhvIJ
oLeZnpq4i6k1hh9OEQ0XocOwCwBh7DwXuUZTig6xbj1zq2hKZwbtqnVaYjuJe/DH
EsjwyXpjHcrY94yjIrWfiMRrG/dUjt7bBd3iPSvQKmZVpAq/orEg/l2LCREyabpt
T0AV6YEw9b8rU5PdOWQ28wCUomRtrc+oyulXBICjKi21UwxpTFi8q/Dt8/VcMybk
mxQemnlWSyG11IdQnf9kSK2qAtp4ah5hN6aunhmfIxFrW61Brfk0bnYIppZ9lR6C
f/gVz3BW8HstNpfbAzKetHuEWic20Iefi7T+8Z2OkBosgY4gKSWLcABCmFVLQKAN
BVe4GsoERUBneQBDuZfPDtZXIk//U8QgubS10sMmz9K4sw7woa/iVacxMPZA+S1l
DMhYVe9LSc/xoAxdvjAKVzvUUlMsxNoaezEKYiO+CyemxpGt1LkKw5wWCRHVkk+I
XLATPLNkUA4UN/9keuje+euoXXJxitO7NH1wwOy5GY0DU3uvkjPdvM9+dychU9eO
aYsuvCXTjOVha0S76mWMLY+iRqjWgWztyJycBVr7P14f4A3PBUvaPjj8DdK1rbBQ
WfaiQj8RGuICinw/x57MoKlHXDcE+3aR3YjYzTPneIomjNRsm9uNOAqVZO6MojC/
U8RFiD+FRP5X6A8MR3xpyJiu2Ag+pz+XJH2lXV2HtNZMG30oV73BRPCofmcosLqq
qor2//U/0I3m0KRMVJPUJe2tK/I3EUXf2jKJhz9MwOoql/EuBljLXZ5w+U6JQ/31
kx0jYStZ7T0joXri7o1kpvxM4kj2KFbPmpZOrv4tQcDcvXlymxOX1KXrnrRyJlZU
kQhhF+QIsvkHwfiKmtvuCwfHiS5XvBEb63tRPBV5kKcxJu/3MweIliydtwMZh96k
vAfDFlCgWhbnpZjzZFpHJN3dhu97PvrVf9lczu2dEHs39YaE66Ss/GmiPeSRIHMw
WHQmkwjIkJBMdYZU3mHv4XwVaamTaYJosbmZh5M1Cx82Lvh3rgJOtuXnm2tGSZ98
RHOi0so9K3F5hKdPdWULCuzbe1kMx5fuUpQUFzl9lxmZWtuBxXN/+P4MwQvSSfj6
MBQirkxvDSSP/4U7LlqIwQDG2o8ZkcDnEQHxGNlJ5HxWTUZkacRh09iXiF+GcXV2
rhWZZMF8nYrdGFzMniOAlLWRzXDfgakRREWRg/RX429XehKAi47KpWxQbE61NivN
VHktTXHAp65XIDUNCibRkZwle3USZ70o8TSrKuMZjp/IXWIyJEw5+RISsItSVxZs
VWbIsW/qc0DCwwIKi3brkiAmdCcEmJWttt+Gjjc/dWZ2e6bEtrncApra5lUmEer8
O7JAAs1FYeFRQcBDrzP8NZNYe2759kuPe/jOJCo4nMVdc2funDeIbSJO59DApz+f
4Ak+wgO9X0Ny+NOhuOdxUTe/vJfXcS6jhCxkdIvicndoJdznU5ONVZ+1i2pZLm6O
N4HFvIdX5rcgxJ119qx+RjUkGpC1WiDd+wdlc5Wb7aF9YaqB2tZqNwvBY3W4SzUQ
/qX/Ugof157fjw8xVSnp7SIeXFdZPBsbqRl1a+mt9axSC06RvM0rR+ZdcLdOYulj
YM3lFuZadLYeD/jxNRY5Kn388rZrkTpRTcxROyV7oqRdgsFzR4ilkh2a3NA+ECdy
3JYfQALme/EvY6fUiuySYolY4OziIZ/zviTQ/iYbCVQ8WFOjy7AljLjWKqV4SqlJ
kAHzXVz8Wieb41AV7FYfwRXr/KdXb/XDZfsHiT20klRMXv25tV0dxWxWIu3iXIkm
M/S7FWSfwCKD7D8Y2UZBS56CKFYGFa7WRbVO/yZkrSkJv2Z38nShsU78yiSqxebp
HuzwcB5IEpwglkNjped4hdPKoWpg03cD/Tibm0WGfkAtlzfBL6Nb9xc9BYSAHjij
0ntr+4C5sWrQsVL5AczIdRimAMX8JXYXZCNOCGA6GGYlBAG8lOVfkr/KeLJxhSdy
0os6ZY3MOGeQVTPyuNnGcscurCp/O+O3NAtpqMeSroYTpF4g9tSSimqRgfjV0EcB
EuSTXML/Hdn55U/SNL2652KSI3H8TuUc7jN2QycY4KUQwfOfOhoKDH/at/HVG4Ch
J9lxe9d8AEXcu59dPX+SIWxxM7NidOvFVBqbrZxzBaksESr9cgfapPak/6byzBw/
Tyi2XpqFtZr6P5w7HKgHRJiVBmrEtHV7Y47MApJHJq55qggRMedZEMCvbOTaPKCG
9/Z2oOMg7WXj7VmdjHm5+y33KUVxA/X56vu08x6tSHYgvmaR5xd9jJ+2mxs03gF1
2ZZwAFmjHXlSXuwId/pFDuIGLQFFDk5Bsg+DHiRu6oTgOGtA7pIaxVwIrnJjWN8S
/2jKt7zRxxS2zqOnMRt3urEOQJaIJU2wITyvJXrdt/bW+i+cu+EgnqP+31Rl1Iz9
5wCcEQDVcwRHSjPCxkWRwms5xB9vtz9KgV2Vkgz5Cw6j3xtkhdHMTlO5hIeAZJ0b
1sTGhAOdqai9L15sSJp7ZWvzWHah4U+udQFrzoToadsMr6Et7ZbsDfWx0MF+2jAh
7715YLPEDmI/BUExKb94tG8fJd/IUsqO//NQEhhCAehUYR6gX55grpHmIO57JSRw
apLo5hvQ3sU/3QgGqSvaLSkmNhxTuPgbx5nPZwa0C61EIQ/aRIIrIWCppsEpCBLj
ax6LumUfmP6yAxNfU/LszxiguAzF+XfGFjqwyv6pweMoiUQu2B/WcwNhZjHSJC7k
pBWXGT2CBBCwd5KMCBpTwALC2LRi7ZSEL8WzX85svJARBaNS9jgPGdqiSKCBvgcd
7vDTygxj6CgvF5WalIcgtkddqgHZbR2gcmsLgt060HlYIwXXLv158GWv3IkyqUlP
rCCJWDnmozvV7P6zDMiv9axEJRirRM/BlgIlJtGE4vGmQOr94JzyFYj/wIq72+4H
Kf0y2ZG6KMQYZm7ALJSdmt7vukT+H8WPL0d7MofoGkq8oVHeo/uRoocvmevu9SzD
hjSDdEKbZmUnunoseqLbk5x0WRhthoyrH1015cZyenI7SC+2ZgXMBAMchN0i7a6J
VcYk4Hi80HfFABh6kicIp0cMUIC0ZMeVuvjW/kIL4fc+GO1ia8kBhGxAchvGF32W
b+ll7tdayhyI90O+Dvn3iAVVREFo1MM/wq2OiXMibmIy5jy8S8b5WiLhj9CH6+zB
wclhJTCwvMK2mee8uipa5KdNtiRd+DHlpjqJWNDW8Yz/C1mmjqd9vgx/66qM+Wri
zQOmminEL7Xjm5pwEO31iIQPyChxdnzgLoQhFuxpv+uJ5AKsRy2ewhXG736yzGAH
5DFirAxD76xjzSs+BpCptJc8YW5PnfKG0a6VC3CNc+p1Xgfe/KZQTt2srE7BWx7d
8kCf0L1ZQjbYbrt1R9ENjGjymUKL48z8e6IZJxQkgYvBhqDLWq3vHWaDHJhh+GfH
IyWWW3QrgniOqMA5bLdzKd1YXRzAE8f2qLCxCPtLJ9t5ECL60iInouIT9/V2lPma
H4rHOWzfYVjjUz82xoDHjQOYOPjH6bL5ntisOQPetrPA9pj93cJ51UQyKxKhj1c7
auQt48QflnAAZGfqykvfUfNcNmoxJM9fz7xr60KLG/eTp4/BiY+KAU+dd/O1+bn9
O2Qk6tjplklY3jwr1RgEYVTtTfHjkE3nF9zUJSVmoqaTCz69NWbI3TYQMYbog2yn
B4QkjnVS5sPuLD02A0REbeVHVV+ck/aM/mIL5pxojzFwHGRH22eIsr8pskmA1ISZ
oea/xHd4o7uLpdN+E5zp+pI8XbcMyABTxm2cFf5s8BN7EoieetkEEhvpInbF8aGM
NfgqwU/qNXA+sMTiQO0ESAwbGYAC6awFydvpBJkOSbMeyvLAqBdhbAIY19AG/REH
/eCDq4axcpa9tUhBOXtzmxQCixTRgNJYRCEMC/o4L0v7XMdyYwQM7mAZfZknVtDH
2HqgLBhrcdQ7f7T5I31QgTeFNpzi/TGjckiwN0J5tOSaxBNd6hpsWDQkNxEZx98i
Cdj8rAQiBSUs5gb+98/OKNl2MYYH3LEw789lFpbi21wN3Qk2i6phIB1yTsnHmTWU
OCZmqSib+CjdX2j0NLX59lKBmY0cA/Z5RZUfDgDYHE3hP9QdGU9/hyv7JoZ++1rP
YcbzEDWHhMhCo35BjeobRI1qQNVxaAp0yBBywinOy9vp91OKPnTW3/9NbltX+pX2
HipZ1DimxGS2XfzD3f+jaCUJVWHtFKlKGiu7y47o/WKxaznjebR/CY+nvVU5F7P8
Rh0VBVfMnNOob1oFYKCRgy6JEBJ0VEoUNhl1Jdx6GnAsfQIxC+RbdNFt1BDQTQo8
Vs4oJcLOwKVEsRYgZOgjVBZJWJSSU24eqsbm8AFLy7A3Xt2rDz5uCiLxLs8TCCrt
EYdN+mqFuBPNkZi4Zh1GEoMyU1c8AuS4IcjoUk36b+6jrXqDjg8Q7n612oh6Tth+
GBT0XpKqgtgAErbBVt74O0b4OgoYKgbrH5dKK1bo0aORwi8gQgJUAu38kk/0vD8P
7QywsLc6OdVaPWQK09HlJesh8Z45JRxbVLXtT1Co6mk3xMGqSTfUWbYBWGJU+jlL
pyPfuNhMccl2hloMdQTiv+ghN7FOeldKiZksLK/IOBVyOTL/40gYgn0gko0vXjtv
3UXLd/K0UACFrI94+j0ltHtp6rRFotdgV9TQYLGSCZDFyckdx2llHWE42fcX6p2D
xaGBwAPz1qM+aPOSfA5rfHBDrLRD1TNyvSObRIaCl/HmIYaGigrfCAVu4b3Eq7Ud
eybP1oTB5q2W1sTYT678n071BRs4ZZUZbJpVZ4FnbB+FucsfiWNUA6fbLEAqBofd
QBSHTIP1qIwzBRLoOOJd//kDpIyBmx+AiqNvBD6yI/wx8LUjWWGS1oa1hg0zZ86m
rT+jRSBzsHQ4MM1ORTaKEitv0GjlYinfmKmF7ar0K/IH62FP2aWIjx79u5mnCxLn
mPTdcN1dVQ6sO+d0caV+VVzB62RoHGx+/zfDh5Rhfk0nuqe8+EH76HExJ5jgIB+N
NMoMSqQhnnm6OGI13bw6fcJCtuuudZclAXvxbF3QeIw1/QLL7sbjeW377GTSczEm
S9oSI3QXhTHQZKV6fDKs/XYmdwVeql4ftL5QWOEiZHt4JpVhGhfDvJm6eqAixQ/P
CkX+fLc1Y2hUuhnjH/z3MabH+iX4hsdDefbA2EvyQ5+rf+Fciy6FLqVd/MGKtNJR
aOdsVSnWdZKinO3xMFaXPRncewhPeXMNnMb1f6M1YsE2vXz44EbWjMo2G1H8KsSO
EYapV3xJgw9k/nQwO4MI0QGBiF2WsOFXxGn5nPUJZTb6RnaYZQwxvDCsKNgfeEZl
vmDEwIuZ80ehF3A2ON7suEDH7HMAiskWcLXULFSSAuhM+gloWYvYPSqOcu0qtmw+
MmnHDeEWnt9yOxi3WUQxBOB77mPqYoOpYtrMqDSC51HhQTA4pfwOReR5IosYa2/+
r1qO0VEJjlhFTSWEUDyEUA3jfFshdEmSSvqkFaHlQF75cZRcM/CIYoydUbCiogW/
0iq0XC8BRij8iKiWA8ZsyOe8LcxKIifP415s9bp3tMzDHTcEj4Q37ZHpMti4vm5m
CXfqijoMkJnirzVDK64hVxMJBghAJDk/PP6ureKux4LGXO6aKS7B+bikzgGOh83+
d3+QxIln8nyExdoUVAa01rI989BlDgcgvB9n++6xzOj3Bl2eyU9F2n59dVO5MskJ
vU7ilTmFT1drjD3W3VGZ8nDC4d7ZS4VVwwYBwWH3DcJqinW4P1t7Ygm+WHSE1kHl
Lbdumhn9pJ8f6Wc2Qx4BYGxTlcCV4k/CCxFwNzh8l/eVa8QtnxsCmUwuoYsg8nsK
hpgqKphDbOAl5tlM6ZzhoWwJcc9OFvr4VZcWvBN8yIeLfjlOgCnbleXYxxg4atLv
rBqaaFPuVa2CkxIAML+kEYWi8czzoRgYSvbd/c/a6twBeEtSYVA14Z706GWqGFal
3Dk7kj4rJDi3wdOM/9ZETy4wax/r+izkfWH7U1GCHTAskuTOoE0DLLvD0sG1x6hP
IIynfY9tSgIiPD8n9yzmtvJGOxt/Wl2lMnCgP+p6j/GQB8DG2bETyS05LYY2attz
u/JX7cYEQ2KRqnGLjKSG7atGYFoaIX3UNGBK3dYFAPSnsWquQ1sBTqcitruM3k15
PSInLlz2TQCwKoJ8N+NOSGTjJpL2YVREDyV1t2gGGIm3lD4aGvAEvpLKdlj2vJZY
ibgFRaFSxVPZQ5JuSf9v3foIogZs2ApWHdJOeop3+RcKuGcF7KP/o6f6Cc7oUO1N
VQMBFFJlkpEWLotPHImhOO8nabsUr/BSKI+MNTbpIrqFXfGdMoTb78hP52GuF2h/
DiKzshXJnaJZ3lrvxzQKNH6moGl6FTwnKxSskHuq4FPdM6Oo85BcmSR0OkU8VYe5
MjZqP53S6ABZsdVKdSzDDO4ND9ojprHACoCWmrGzPqrbfeeKsKXKA3nZ2ayq7AvV
pYbAP4/azOsZxxyE0TGdQY5NrBu43RMOaxP+Xww/DhlytEnOvEou+QIb6d+6T5TY
Deoe3epnCJwMDiBNXvse/mGQ11QtP5HwurE7mdw5n8MvXWl7RFXbvEQbAHEnshhR
BopUMN+85Z8PQMw3B8QRLF0yLJ6Qp9lbLBDNY88M8RM3watV4fO7UfgUH1eXAnXt
f0soHdj6H2BFqy9hUYZqiMIwt9wYwkxs5qO9gdE/t0lOzzh6XxxefjkJXdFJBdlb
M334BhkZirH7F4PYSGj5kWbJl6S3W1Dc3/n6sOxFH/bCZ8fb15/4slYgRUvS/YgC
q/PDuAYzrzZ5xUf+GSFgHFANt232lGd7Zkzaz26OHHixa1xMSpKOm3YEg5M5Pg47
3nYs8mP5eoC/6BipM00NpZTltWQ9NuUM1W191MR3DIS6ckbd9SfaGWHs6LWobZQ6
sEyYCTriJsYMqWy4WdO0Gq1rXHovrPhd7EPe2BIdKn3JACmB4FzlzJz8zEJaUVLl
U0rVQrBXwqvGnTla80+ipI/MEm6jgXxeoY2S32zUBT/2RR399El6CL10N32eLp/2
x1E/cWPM11f9nqt8Lhp9adUlcop2MOfnU1/v0rQEEDabK1AVyrfJOL+LmMqg5V7B
WPdZkOF5DVGtprs97N7BX59w2/MZI7Bf/NzM+mvHWoIdkgV8J3iCLvt9I6GRIPoV
AQDObU6g99JrKNEg4vI5DVdmSzWT2Jutl5EML6HPX1fvgO7NvWFlRwmv9rg36xgc
UJUyIhiEH2ADiFV3xRKVfqDxHSGxpe6icgCfjRVTEQH6NND7HpcCy7/6TGRYz/K3
lVseOYFhfT9BwdqPwReZZo96gSqQKUOAitC0Z0052Vd//mKnaMzGR7AWdoPU4I2R
wgqjnte5XtWCUK941SSd/TIe9wFM27nDLhDA4GBGrwX2pKUUbD+TZ7irEPxoILVb
+DXyFwae1v+oM9olcEPf6Gu6RVEQcBz+gBXUy6oDd5Smixka5Vdm9+NIo891Mohm
a8F/mvdDFhxvUYhJKQW9Y55BfI7i+4PJ5hPGPVHcOh0NfXNvxCM4rx8pmQKoSugv
erFU7K79/OuqqC/FyBfLuotZfheZclJr8OwiQDaC1EZWcFzXQHIQ47GL0AFIXfwc
TMNVozrNKtFbR6deLZY2LkBiXLMdk2dudwpNS55hkOWB1FNXfM/7E8pZm83mrku6
txM1BfF+vBeDWZEjZmYnoc0KlFEmKCrdh5P7GMJG8eR5kwSjsZNyJIujr2Lczc3h
dsIIRvIDreAZNMLdPJPRQSDxxBe508s3XYd7b12MwTB/YhJIdicu+cyQQ163sFz4
x/UPLx+6W20qN7ezZ5YQrmXOh1HiPXFiB3kzsDtPb0N/DV4tnB9D+aYmBrLPc2yX
aX/Pzlx8+WzUuts/HuHp/27EmVCgh4uoBuhMaTOi0FMzoVSby0zKyuxx+TaVTRzE
UuZjNetQ/R0CyR6wQEEvEegGOKv1xVAzUmfjTPdndV5ZzYKArotMZdvpENJEfTVq
kZdNpzUY8rsmLWjYtxmkDIXCfZUUo3v6ETxM9rWBa50wGiJkdncnJ3NBQDsvqVKq
P9JGGJ/LKXJizrKZ2SLZ79hD3YfnhxdfzSZ3a9fyvGwdrRJNalwyGnsMyJ2qZpQx
7SJ08BlwfWdfL3tzgsUWohJ6fL/FXin8sV6PSDohXaQDrKxcvyqqSJBdhSW+GifN
q5ktjsxjDwiQRGmtkgu9BPfPHFQ3EWtmzOHLoH/fJa03UrG0s+TXw690lniGapmS
3B4JEFyZ4nlZyWiu9pRU6TUYLmP+Dr2AiN7Hu50ictcLHBW22EBRhrer0l/kOg3Q
d/KOdQCBV1R7o3OFfmBapLe/crBIOHhmv3pKxAf/8y47XLjuZIzCsvCzfKbHq1tZ
TCdOujMJCDAaQjIVEuINNmpNlLmm/rozNrdqI9ihm2aYCw2bI1ZxerCPxqf9C2eW
rVKrDHPWXDcLL7CZDDE2ICrwTLUg/uA1o+PNqtkSdwTWGLuhPaWzjl7TtqqTfps/
XAQFlMk5fLf4g+hY0phc8o2rN3qi7+JDRaeQzNbZpdi4VKIcc21kwRqxij9JnwJ+
im3kdoRMSVxkDxyZM8kYTe5dBh650gAi8mhCPYSHpkLV5KufFhvSarpLDSQmC5Su
ZYBZmEOXc5L/aznZxOnFHdEDhVRsMv1QoxIWzNf7wzhRaZCR+GDb5Z3hjo1Q10jr
dk9eVNugK/CPXFunjAFoQeuZEjnbZ9Zm7MAn6UEhB9xxX5u7z/yxrx3F6EsCjy+c
EFAjggeXH2a+/X9JmvG2l+YP6lgf3GC9y9NgnLn6MHLFtWNxPTmdx1fmUS0QNn01
xyMjtx12lGW2kXNj7q1Sx/kUTXJmmpS0TCMiFYl5ofLcFlaeUb9mIlbfw2C7be4s
0OgfcciT/j2E8WhBpY9K2MHbiwX9fLXs1Mr2WNjlklCBa4cD7fZkYpPm9P/eSf23
fRDd3jEvTDOHYMadNKNxz3GK9b0Cb55JSd5ni3Wkn83Hfsl2u91Yo5BcglVDFALs
Ji/rtMKo027UVCdwoedzEgmsePBPR9LG7I/CA3KFMyZteNWz5i2P0EE0fkATqPRv
i0p7QF0UPRzTbH+Dzd0Dt+ZaRtITpJw9WeZ6IjhUYUDqlLmP/m8c+W3l84IkVnl9
/5oDlOL4auWQMieb5jIkyWKmsTHq3QLjcqymhkrvEmuJx7NGbfHXPhAqqjDAF8Oc
geT9Kuw5GtHzoTg+OFY+/DaHbo4HPaUJkDmK+aHbh1wg7GoULxxEAPNzpZejdn0K
QoXTSIfWKsrw5iK5z3sPl2Tx6MbCjCiuT7y+sFOvi7crH2y+94vpa3Hu8LEJFAPj
YOyAhEF3Xr9Qk7xSKONmSjARqHhHCzYcLsZugF6boLVkbGZ0+F/7AQD3J4pK+DAe
BfYENSy64+YBZTy9/rfc5qep/jbRIPDSaABZfbOiD9phf+wU4BDYiafbpLy4nB1t
dhjcxdKV5pVFadh5Xfj7En7tr63z6bfVSZ95xtKv0nM1swQ+xQA9Tlx6p+8jJlTu
jtJna1jS3qXUuXf1XN9dmfBlfXFnyCEordUB4yu66vpV/ZgnxLsx+T3rXMPLS9bv
puIEDOphl5td/jAxMil17D+EjrZD/STqCtD8yF8Gu/2Q7rbCERA+MZnZjBrS+XQ5
lKlN5LxgVDVz1DiDXrbRJ0DHpJTa23NoMUnSnCIN9OcAjIAKAax2jbyhg+TOurdz
0QlEzpWVoQngNd0hjy8YUA3WNAUYf6976TtFb7wmuy/e3o5ExKWsCjw4X0Icla99
YGzRQQeLqz7xPJrVloAJf1p+VYlA5tfZHHYI+LMz5GqYGkFERSx3zvqncNVc4xZZ
Wdvh5OYjJs7i6LlkuPXs8Jd/T59/HG4M3PmZye24ETK0f9GOfZrcskz6XX/pkPeb
Os+7Hei/NDXF1lMbuH5eaHfEetgLJAThD+3tKQYkiDRs8xzieKTGdMnxFI3XQIob
6uw3OrBTKlMfoWcxhZZh4Cq5WTF7tox8sqX6bZp6dWfB+zssue+4WyHs+FSyD8j+
mo2o0Jkfj9bTaDftg0ng9l0kCO1yF11+Jz1iH2GVttTdtLhs005v8k2/ok2ijxHU
jBj8S9OzRV+ZUWzdWyNeoMq7WmCH4Y3z74EeIVdL8R4uxaLPV+OHS9Llqw6/ty8m
3G5121LWR57KprPn9Gy+B99cm7x8++yIrRI7NKa8ZXIFXu/sQkG1x7+P0XZyCJL0
QXV61agKc/e/Fvr3id1Xi7+UgkFVg+IK0hUODdYHEYQ8SpWP97pBEsFR95YNNYmh
I7GJBdRW8uTJwpeH7Jy9ZLZ8dn6vkua9PfT2WkkgFkVZDbRTewX+wRvk+B4Whnj+
/OxLJ0ETPxHnqMvCCI3y9zZ/UMGdFD9n9bw/wOqQ8+POwCuY9SEs+xvQFX3fuG5T
hyxwV1bA0KnPWqtEkjwQx11nbXqQBOFCB4l6oU4V6ikBL1cCOq3R3XyJGZXNkYii
yeZtjPZmJ0c5IRazoS8Jlhv+6g5zDWUIJt4TzmBE/5ElGZoEvKya9gLfQeh8WPDG
Mtjroyrq6MgfOcuMiUf14tWAfy6QSY91gQl6WyqOnRJNtmg2gqn7RFNAJNaOLMlK
ticAxsNQ4aWK9GZO0CRb5WszKzdM/IRXnHEX/xRLeXIEkGD7f/MkBHntCFfz7yam
YmCp076IcKTbZjH9IK3gkwAV2OInJnAMnTcFWhOfhjwTkjY/DphAj6QWgERPsKWJ
Okz3eJPlxr/UzzjUUZKlLV5jSyjPwt7g5c+gWzj+LRxegZdvBYNZThwP0dYxzKOo
UUgsZuk8mXduqmG5LSqqgWLPgs+l9iHKL4h/gKoTd5hvLH2/10N/9xlvXOrZU565
bPspNlRsKW7QimpBspn30q+bc7PHRRckeSWgiI/Kq/b0KxCgWDjz5Z/oIxo/pjtk
MoncmHhujv91gPqN2oueUONX1O0coS9O8qRZEzY+b/FxKMDdyhRJOO95eATW3ful
PbgFTbDKCc7zxu0p5jMaDy7MWTeu51Z9G90KifOW2vUhf0RKOlwWL9g+C8Ffgsdc
KfqidU+Rahq5pmmkPAQDamy90R6OPPI+BEsyUyTU7XqLGRn9mt1tJo2Ak9MRAwmg
uYZOcNMUhMQCOvY7iZg5/Zrhw5+2PXH2CIXe5TJDr8dq9wVQRrmyNPGJdE/QthmC
U5/33iYotsvsBnbMDUwJOo4r8HKEhJIJMMKvdUlRvkZgkmGwe+IB0uZj6UQW35id
vqDIcTMQ2AVtoH/NC9CxhR4d/uUFhRu0jsHIhDEGBGsYKt+LDOxJK4PxXwmGEQR6
SdCkBb/8GQSIb1hjsyvYd6MauvE6IkQ0qlS7o5JAPP/TsGGBsyr6XlXfSWlEfBhx
wj4+6XiyXfYYDGuLg2TB5ES0S3XYW0qBguVS0yKbGxIL/oqVeVW5Wnu59bekYJ7/
lp5Sgw1DJIiDe44VTV3Ipr5TizKLLWMVr3JA/mDv3ekP1tkxoN9+AABdQpcmLIls
SZpfnXU9XS2wMGPz1CPHkUpNFEVrDbve6s0R1L5bdvSvwiieAUJgmiNVqjfNmay8
hvuLM5CyCYfHnIwWFQk72fob7bMDrcmioumHHii5YmLWcaSL2gBAiwdoOKQL532c
a/88KK9pg5o6Qhul7G8IJitUAEKWt/poetWW/PrM8SWN501y4bzD9lU4iboxTE/3
h5Cqj+Y73glUvELFaysDrF0zDgzYJ5S0NZNxZUPXWF6tvxsEJkJFNrhN0JVAkDjz
CornM+izAx6rjGz/MPm884+YCK4bi3wct89nAfCkdCsCqq9VDUl3i2RAAYbh3asK
i7yBwnh311zx3CZ5efoDEelMqbkR+z81iYQXuxRfnkI08IvoRLZJSAyqLofiU5ZL
nVCB9i3W4I+GD7VDinUn7hTIdGCmZYcALIsTRhlkfxL/btU4Y38nkp9CEorupGR6
bvZLXxmlgGEfPP9pcvr/Oi2bC7gLINIKe4RC3nNKiV0grRL0LWUrNBw9l2sL37Wo
cY0AJAJwDyMRn9ugjhjqfMmei/sTnyu+1fdrt2HrzuFE3PVpFzSmeyhxGWpc5iNk
hQB8by0VXK/bAJ1QCgmcHC43+mGCjDGWFE4b8UnJCDG4s9ejE023qzun12l3h4fj
8IXsfRTIuge/S8UWz3Ktvhchd1OHi8xVVvN6M7W7Du4bsNg3VKasPZK/CISnhHDB
8nOSRYdeSqAsMQNCjm+aYrc67bZo347qpYETIBSVSvThRiMOWGEVm1Yv+Husd/Xu
EEaRmToUyr0oJnynD6YDcFz7mXBxJ4mccihm9sJUFM2i8lkD4qdkeMNvUbGnUyho
AEBbwfBgrgQROOL/1B9ABgPxB5GYzrkUGm40xLQ6j1DLI4SFFYw2+i6ijmvwngbx
auGH+iFLEum+e+/g0mlgTAThjmvCrl66Nlu9TMtRtqByvyySyUHQGlBrsNYnPL1t
ZzDSww+tXGLj8cKKkVGYF4y68flapG2PGq4t5vttvDcr3r5CwAHPBhOHI7X2EGfn
TG8tLjGRuBnNOppPUqcG4KdOAKKGjTAna3KVlgj3a5hZoMKOJ4GB7M1A91m8pNbc
w9SKGIHDpLpp40XqOot7fz+j9xkr8awPZOw8mrrV/6cVtJU276z2Y4vesQLMDIR9
YN99Er5tzVHVDpIiNE8aWV959L92z+FuONhVDd4C+CnQ1ZjdL/JObTHXKQ2vO9c/
JOLDDagYpqSMthqXGPUz6M3CptYD0jmha6E4XdbVoOJobs20aOrxriYWcuCxr9DZ
m9GqaieWGy1SvaU9zY0fNuAV3Otq/Wiy/huEoQJe8pYnoZrP3lBkU356SaoBH1GJ
QSnoByoKlcEmRr46eh/lFTN4YC7n1e8NeNsD18DlPJ9RlI2An3o26bpmIOcBz0iI
hc5GvXjHmepSEHuFm0DegZhsTNJH1m/TBewysvi7Z3itzFxktgkPN6LJ6O7v4mBH
M1fkq7uEFQjMw65TpwscCoopXnSA6NpMAAHe7cJbTFSZEpnUzWZVP1EdhlAA9gt4
qc5zcVljytqlnl0imSNJc1Q/yrhEZdLaZmrUJh2A23m+h5ESlTbpV/7EeznZn8qx
TzblT9m6mHXCCSEOVTPOXIeqrnOG+iBbXwQbMwl7N7mwD5YgazN1NT5N1Qq1elGs
xxM9Y/ENEs4ur2UXS+vs9B7z65XzE79RhIqfzttDyndsFdWT0PdLlMahrcQZRDoF
v4kom7jbVmC7mgmznTblV3WtLu4W+6ijJMp2RxQHyp/MXu2uYUCTJf/vjfqXln9K
lRyyqCSNULYLC9/O4D7GXdRB7VIOVNKFIZxu3z8ykFGJYYVno+2T5LADpPGwIVxl
9uHJEOLhIB+ZygWgfM/Nq/uMQpx2WGi+y/WXoVJ77sputQnfbBw6hHXZ28VvpjzJ
ZNlgnlT0oxj3B+g8E9+YTzc+x2f1a545WHRUPTYtoxDjyOdcpg+lh3ry1g3qT76W
YJb15Ab1YP/G/nqqcNbEdWU6p7afpwjwEnfdKYBIDhJR5efYxY3zXBUTkJ9Avvsg
jrjABUW8IIohbS2yBLM839/IYU6+wVibAsAzSHvEtRxSw6f16dAKQfsZ5rXLKMv1
39WnM9YsLl06+5t6REP9DULvT+UsnUIeW5M4uhgbPj3GG9nmL/9qH/5uMbFqL4su
WJvZGF2LQDZ78P2SxLJiBSwoiDYGAwoTPasOFDFyHMUrl/Xs6hJRGuqc8OUKp4x1
j+DJ2bsUsULt30W7la5P6yiLseSFdumBM4W6jywtX95MwZRF7Fe9RADXLbUCghLV
UyTrrz4/2klS7HFu90mT5RsIPRl8FVFCIAFQwv71y5GbMyrQHtuTbzW5Lust3Vy/
L7MLmD3StgD51WSpgNoawq1jM23Awkvss80FWwwjvBAoAX+LHWXDtF1VNOQumhhS
3dnoCCVRRBaN9XrMbWokK2L8IKh4Rxhy1wxVRM+4UqPGQephp0PoVXUuzD0GKF6J
rdqffChmf0El8va8X5zUBvSwNyv2L/bkchojjBWljOaRwOwWJTTYfvxYDgA+b1l/
FhUZ5DaZQPVUkWBlXX935belZHzWhyr0XFbyA77/xtpzTMGv5zoj+0v5MuDRIJUh
jR5V4dAuDgWt7vrY38ZbZpAHrm/6YcxWgSEm+zBumj9uRMJu/sfJoZiJNRaKU1/A
andTPsADYiGUo1dRi9M2lh/MWWhuqJqvTVba/icyo/fmNdc3MrGUcN6DMXWxaTYF
ES4ohRc/mUvefMqnYuY6D5CcxnvLmS0w4FM4q+BMTcNlJVzNSXloEKkI9N5z1XOk
QnMheJWOh18D0pBrpcKPy873zENooHMFij5pcotwqIAhuCNoOm0lqxwfKIldQtXw
Wv8pLNIHjGejPSEYenlQcQsQRmCSp0zjZH6TcolIAv6otFBpu6/LC/eaVX6auw6A
5me1V2vWCRFFW5N47AgXFORslLxkLCcOHceM3dfWDdn5E1gtluWhAeNrHdlO8QQv
PkFDdcRIsS94V2k9SNcEtdLlhXBXVlHfpDCCVTKNfP5tBW0Vtd2TbZ+AJ0UjL4ef
Po9OGMC0mxy19kAum6XEFAbKkRCnnM7RB5AkcoEiM/m57A0hcy4JUrkBPaPm7LmM
abcRVbMjzR/5Q3q0s9FyZdFVpKevJ5B7Z79Z2Hh+OwgfWJ9yywGF5DBguggjoydI
ajA2Orm9fci0X8OkV9jvtXlQlbQpSXMnkMix2lThxsLArswTIMuea0zyIXiXYXUn
hHBTvGHrUSUlyU1WJKBCeAT8ad8vIYzxFm2cKKSfP0DzwEBJXvcAb71tGmn1zB+Y
kxcDFs7ual+0X/2uLwL5ctIf2h/2YALy9Xk9VjMbo7wkI3Nfbl9h50TlOzGkwhiS
O15QzuMHLdT9pwjv59IgNjcloos8nzPsCQmRifH5hMMCfc4Gjaa3hkICMtNUn5jQ
FGtgd9fb0TCEViLHpk1SO3rIuouVy759BZLuiOYGybXJyHVWqVh76mp1ZxTSfjZH
rW99MAFENm+82Fe6WU1Z+tckBHd61SLFFH2K5aCnh1iRqC4pA35RTWVoX2NIx0r2
0+QPDXhnECQwtcAfGrPCbaZr0Sw1DWTn5ZbXYOjeKfpSEDxjY0Bu/QRDqsDiGqe3
bh2N3ghChalBzLbwK3DF+I4i0Nbtw4hictWis72k8TUL37eNuqiCwvqvXH8+83D9
uSZ9tjOQvvEitZOhFtQDL6PtyT1h5mi+vH/K8S/dc7B5FgkSz64DVMNQMhmIP4Po
ELBAoq0xZ+lXskzvGNQSThp1F0pW8j3AWasBZ8iETKV4rs78AjHnQrRQkz05Fe51
MU+MoBfPLIyzIw6z5qYoa8qw8dwJImjjkNdErOBSOsUdptS6VQTczTB2RDJaX1Ym
kpG8KTmixFdaIknwgcIwShhDGi5PjLk5gnPt6mQNMjU5XdjsAYnISvmr23ZNzoBB
eHMrpJ9YpE3ow3qVCDkyoi0qLAb3evaNc8atjaraXLvaE9uny7G+SRx+jtms2Z/p
th4eP6aZ0VPQ6IBAZeN1RO9kkOuHr1JyrgUC0mk8pW71A4e8cxDHzhdm4HUXettw
cFzQcYrlAMfDELMQ9OHB/6Y3p6gaPHT8dAYYAI0OzISpbPSMCjvuFkBgwMTrrx8l
O5kGrbbPYmQV0aiPftpFjCK3RXNSFQy6xnPO5CoODhyr6tNld3q5GQWVJS4gjdJk
BShQNOA1aDgZdnWWMzNTwJScHgdpC+94xbVJ7LH5XZ4ztPKRVvdTeq+dfgS5KG+N
64Rge7LENsITfg3BlMC9QbWgeEAL5wt5kI7WPJ3/WErKAMjq0eLQJIyzrnt2s3eB
ztBwU/pmzzxpkff7D96Wurmr3wGoQaVZ+bZ6CrqDh8eg3i2wuTijmL6W3WDcT1a3
8du0ZuEy8n0otYmXWpNBYciNfSc1EmM8CnSPjZE7Lp+AN7k0Ye823fdwlTYJjfSd
r/cjXlJCltCOM4U91igukzgb7C5Hu1Q/LGGYB3l9yGiPbybVY5vyRHvKcUKzqJ/v
87YlybfFLjvyzxyCfad/HdN3+Lq9JZJpbI4vjXA1VC1jV5t8DloqJ3pP9qhuCJEa
QIZ9IlMTpbZCwd4ej2L//zyU3t7VdZymcNjwNzQWCqH9UMWVYCLqUlv0/+gc6KsW
I1mhj2V/8z/qFR5dCM+zkQcuvExfHTKaYk+5xYeT8hFQlAdq1AgVmwNR7eCJ9rvu
oCQ2aZbCU5yO6HvTATAOXqCk+7mcs6lpn8luB5bm5s+StSZO9Gs5XW08Cd5jPWXw
AuukbQiTVAOvbT20Br2RoBB264yil9pi0grOJcAdwsVtLJJkc5qXcUQtc7Y2VzqC
8eGHvSJADz0evRKkR/ln1nnDdXEz+kCVpDztAQq2zq0hXKIP2cwOOePAOiYbW2vy
AAaeIYJ82XdnDQrqKMByG3iKiV8tWNvV3A436ZoQREunOTyZoX2jhcK5yoQ6zuQ6
E0+lVi6ujb0i9RMH6BLThqWudubLnK80n7sL4E8aauCYUY0Zfi8ubp526B6vJThO
YBaLwoQIKIQQJoRvCPMPrJeDIB/Q48APWSQyuvKIwVHiltpaj3Ren9T1JrXb8GY4
k9uy7IxPOa8f9+XcrhTOZ43RB/o0reGajGRHyRFVxzIAO0rKwzFU8eGPgEVuCRro
vqk+IFA3jIog+EDCAhaz3K3Fx1Q2EMJzbqbqjhTDXX8rCU1CDiVZkdO1n+FMnT61
zzmQuzcttKUGDxFXaPqokIIgXyUjrAwx8iidTZDyq23wpcAkpDjlxYS5BProptl4
E1H1y44armAhbdSy636IViJFrHC48t6tbeDrBU1qP+ECPi4wTk2P/xrl0Q7JKS+B
T/vT58spU6H3EcSdDAsHTb1TZ7xRG+Cs+ayoGLqoezcJ8zZQG5qJajJilqLli400
6obY8kWzMclNRzQA07j6SK+ht8RWGoMVAGxD10MsgFkPj3pnf7PhQzHkiprjHzpo
Q70ofjPioYNra2SnFMSMUA+yI7LesGSTfrzCLlpilK8pICgFZ7Or45Gslu9yrNbd
aSD/xFrIKJ6h6hDhAD6HwDYe19/pcAWoU7ZQzXHsxsrTCycZKfO8zpHsBUfuz+GF
5hkS6nnLIs88LOdnenUruf451KLwcuKPlGqjkBJw2W8/zWHo6N/Piq77J4rOdkap
sU/y9GlwTTNz5LutWC96UQBdJTx4cU6KjMoMFFZFCjghZb7INy2K0YcWnhkgcazN
3JXrpWCedXdzVqYrLAaKtR2bV5b14Jijotj8v57q/y0xW2gFbBJOz5H31Y3qe45x
BV0T3OWcSprZf5yECN5j8zQurTqHZGuzzxbeV8ekA4EDToXsRdoJQ5QpMtuJNA5N
oqrAZkZ9nFh8or3yjE9BNco94pakXLDFKI9UnlvIwGkQDls4JmN1VSLYolBaTUQi
96y9YL3bHoFri0UzCJqHVt6I9/HEzST4z1Zu/xDmqZ5QE1tti/E2FBUcxc2deSIi
ewuboZ+elDOXyWASQy4x5oKVsmKeP43xnqCKzsdjCYR3rnmRaMVOd1Pg1y1QVHfM
8xciATps/zEv/3ua4k515Pz1E4FBKuOifKKqf8+zm7V6Znw3HSrrfs2f3MIFIs8n
ZbXrwkKGhR+VfSxDmmua0gLIDrEZSxnFxn/rqd4QnPl8oSHaUHc8aW5JmwN0UrGv
4YMZM3GRe8s+bJp2/JkcP1YVn9Is6Z9xFFcwYTT9XZRF6oGH7Y/jG6ldYIztKu4F
JrPGEwP/mgBLxs8Dcwuwd5VHbDGoavBAj1Q3KIQhLzDgaxLY0zHids8V+/slZpH9
82vF+0NEuYy7XeTQJcSaMnuVoDuTDSMZpdnfTVefGhrYPpSs6XRqSpNqAoAb6wzH
IlKKhC15mxHVTAJE3cI1ilrWNYWHFgERolzUu8eGlxAjG2qGWJFqDIMlT9HZdhoe
FyHQRv0SvErtmpx+vopPGpCA2MWs7DeDjR4yEyphctoUHPnZ42nJ5M7iNnFrYnnV
I5evHygD8jHT7wlNDsJnFxNW4UB1ZJoBCjcRaG7qvlYSj9qEVvnugcbNlF9i4ntD
AuLWUwNun0BroaFO25bu5NaRxDgW6m1K8GLXxV7p5YEaJfoOeZ0ViE7SVJZOYLSj
LEZLAzvdy97LsrqI8jhomabBPdskeXDjwO/P9vBm/f3dmBjHM37+BBoZeFMu9KTi
9ZbdmSLPWB1qqUyEtWMJEKPchN9Rg6MoZA4nPV9RKA83VJNMe2uSbQmrmfSr5EHt
rlbQpLLBzMrB/EZhm/JpV01kpLibwQJEAECNXPemJqUcjjNt98l7CxrPaoNWHWDY
AUf/C/F7xJug/p5NVotu1xg6RO8bt+z9yMhn35+U51ENNBcLRVmzoB7qI6WpijKG
Xwy6XpBa8LNAC1C8KjcYBEyA56I4F2qcmn+38S0KK/VFVDM9qQCNKhploZWPU7if
GwYf7l8qYK5eRMY4658RLXyToRPJNC5iJZRXx+SoRWW6i8U2grixt6JtUeRI7AAT
2WvowlO8i5jGPH23mIp0mzhQsgkP0uQOKQfgSsFgMpUJ8sS5ZKVIYGG+hx6j4Qpq
ekJobeFwwjTBB2ULXF1G6qMBRzN/Z5E4X94ACrATez57ES1d29AYKJ04iedl50IE
QNL3Frde41cKK/Erdg1V0MVTnByIoivmCOiW9TIzJA7rSEylWdYKGy4CzgXfEHpY
i4dlotzziNABF06or/3lDcTeloa3FSM+13nvQvsgsZdRx1ksrB8mJurcCZKqYkVF
aL21YZ4Joohh3s9PbXZ9tWjh5PgqgLPAzQaUDBA3G3XTIRE7C8tx8eBCA9xNot8f
Kqm8oZB8GMGc5gIGkPNAVSQiXl3FdoaNShOlAhezlVQdC7EX5Bn7k1XoC4M1VwFj
acaotXRdJcd+wzqHqP7KhDV8MFd/mI2EzS5lAaRJZFte/OiaZVea2FN8mNZHKjLc
U+ZE92cA3FaBVC/kvNpmuVSqoIBld1NknFR0BruwccIRjTqHzkxoamAo33sW5H18
7gvrFnNkaJgfcb+nMwDrybtti2HwKuEqUYJZlMHlGDncULz/3/BrsahTAbTXuaRy
3hqyCTFqQ0qMbfGwPN0lqi6IdidzApJufbfBvnW3EC4c87m+ic7l+uXfCiC+0Lpt
g05KjHNlrKZG9WsvYCrYb9QbgqI/yu2O61flDrA0xq0S1axGEUX5VNizUl57BCFe
1gZNxdssQLkm3IzgXsQP96wPJxKHcUJDUgRUC1LmgKwpSASFooxxwCldDz7QWTVv
1JYqR45+sybetHI6B6RRf/w3HBwdO5wIsYDiU7rsEIpoZAwEKf622KyIL/7QKLO4
7dd3oPUeozQ5eTzGP1smACqhgioMVp7cYHi/K0JTu0qUwJVGytEbJk4OxunP73fb
hedjl5LV8BHr8YoLgp64wNyjZFVoQanfGZOIShFaFq/RKQj2Fr8yZ8UrwdCqWb5p
XqzSs/NVMUFPmNyMR5ZZ0c2x9jenhj9Z9D3uxeq2VCsJSnJFgNLSLT1kHbyCEf2h
eVa/L8tbPqo+DmGZg2PhCItwZr6xajpGmnjMqfpSDUy7sPUoLNfn3lhC+ef3K5nC
G6cR2EW3s9MdrGxyOq5fa+1UXxcY83EndRYO5KjOciPPAMcOJtTlBoM4Q6MgDM8C
Htlzj4DTjfvj3crKwTP3WBWjP66pMQ5kZ21dMzD5bz8BchoyWlcmyZUOQNIj3IA9
3Po26uwsnb5UKpi5RSv0EArf1BxbNVKS694NsO2N01/I/S+cBOGrV+2iNTXEfJiD
X42LKh5lMpL/H2SlGSqcCvv7jgj1CerBJn8x11z+7M443t//c3S3R1ioPta0ZUOc
URZAs14FiIRumx5/RJNMwpPT5l/g+ZRAGjSKfBbgEyRaFSG94sQkfLHHjcPao1fS
E52F071kNdQvSvZ2s1XYy3UbvyQR4la38paYtq94vwRIyOb4LdpvVmrla0GBIfSk
tmYc5+fl/TP6AA5M4DOMsfF5vTduC3ENMkz7Xf8m56msjS6IWGG4ZEwKVmRI46Ob
0tLVbNmjWhxDyVDyUhxn2qsN7gTF89zmhZ3g5cB7XSq7bvjEnjWgIdDsbnO+KbDC
ZCpHauyU1/3fjJBB0e1SUxsnCmgqRXOpO5W3Rgz2/69JXg4waS0wtP/Ps3BLC8fu
7FuSiOX7JukgSgsJ0q5r9rFyiIbUiYBHVx9O2/T01+HvdCxmPLDO6L4cT4tYVl0l
TZnXKy5csjnB6zCTpPmAmclMWkQp7gXbkrRakEb2YI4DTQ0iqo2gft+U6gU34B9Y
3mie4bOogGjjDp/qJqD1VFLruv7VCHxB5xXdKCn4+3yHnU70PXuBTDBG8DfGrPaP
P+A16zpFx1XpTqphxxZjFKX/ukraKn1LhOQjb4aka3NbjCKoIowNwLAk7ZC8u+vS
Id3Pteso7fPHtdtpkKpbHX4D7qSB4Ck+KYUCHeqHGYq4DjW+LSnjvFBBZZUA4bjR
sQyZl9iIpjQbpY/AI3npKPxoyeUE6DWU000oAb+nFhCc1L0DcdkCGtO/G9vNOjxy
rBtXBzRKYSyOLTqU54A/ocmMIoeHAEXeHMlYlKsKOrsTUJ26+Srzl5pQ4VIpvkTy
cY9DQNVPYjkOXdrtbIeLbP6GHD1mnHVU4/zIC8AWCJ553CUlf+m3P4SlprORaZB9
VaXHeMtr/oIwV/XzWOqfBZTrjHgyuNuodeuq1TLU6PN82C8LGEkkfQSc/um2Bc3r
YE5lY0b14gsDOKoG7Jnj5cXTv5L5MQ3N4hdnIlpiAvW7JXuzxcyLDw5VD3NwQWhB
AVQKV7RKHmhaUQtLny0Y3bLCzh8uT/k/hgVMh4VhTwsiQIF98KxLFb1NUBP18e5X
KVBImJ1GPD5Dd2PRsPesCH1TwiStpbykLHFbMC1smgLj93VanxWRfAlFNcSnJnwC
XkaVqufSgpEEYr9m/m+JGu4HuI3gwrEAEhwEfMLjGPpIx7BCGIpT7GIKRZk6pMLD
UqIucd/Uhdyh0M7IBmcYjEOeQcrPhL5Pc9O8q9DldL1USqCM13o94Qbiw9cBIGtp
VTTkjecC5ETfPEWEFVdd7+U61vnL9iQ6dZSIIv2Hl2Rp90C/GGwQmB4WsDbJWlnG
LZG5Olwv1ZspjhTOBY/J6XoxnuFxk8BlX88bVzCm7t6qymGpTA86121sCtqJSVT4
I3JqlVhn2n9kBHw02TfDt2Zh8M9bNhND2ECsZNqhSB4O66ssKIKTD+rAc4keQRgd
BNsSkHOUMkkG9WZEZ++SvX/sVvTQvZO+iBN84GqyrTXErVfqMCzRh3hAJ+Mrd/Lw
Pb0avkB2OtZxDie1UjQWWnX8SZaOXjqyUItz9CfxOWOMKWP7irgA1xifFsvtrziX
T2JT70+bZGlRBzir3AvO/VxBOniOb6Xw/s3now+qrxryex7Zda7jv0d/J0pF5g4D
VjNO446l3oXzKr+fDAx6Qz9H2Uzg8NOdx0NRBTTVLo3tAHbvUhG2+7FxtLuGwY+4
Z2RPOu3BdceMBD5xPqY8zA3OkDbdSTL7yOwqmgyuFEZ0VFqPPp8610VRH4CvMWSF
DPwyjHuNcm116C2CAzxSOn5qmnHVEuLO9IgIw7kbM3Aw61upqdAc4p2gdnR8DFxU
UXBxCnhjdZ8IZhYaH/Nf3PFih9HdaXXkl31tRVKA9CQZXWVhI06eHW4f2r3Pbaqn
I6S7ZXK8M5SgPOZ9OXoHu3pGKq7/3wrmSX1UzH9qTrXD1X/DNSz7MUzQpSxFSNEa
7xxZj18DOedEItP6qWbcFdgp6cCI+On4H1cTGWzsyQz9G72E5poVKMeqmUw/oUwz
SYtd9hXvICHtno+lyUhF3xLVvzOMY7OIzSyDCi1VsiE3e/dzPSq6Xh9e2Vmg+GYI
6SyF0uy9zfO4z0LyTBO/qGUr6HUbL0R6NmnuDCzq5S1TW6PK7pYmuowtp5uYWXvd
dn0PSAFEatVUToNNOEv9orjp+WX89YnhNwIhG3nqmrYJwYMJA35AGJDNG5ID1nhc
JVMAIV8A/1LoO+YHV/eh6zjDK4oMIdaO74LyDMZ6Ml7Z7PbU36OBU80uA5u1Hg8t
nDcvgUk9HiNv8OCl8w1ifpOKOZdA++vJ233N75FdRFmXTb4LQvu2U+LvTQig3Bmy
1/vCANRJA88AjNMhaTg5hSydSP7KJ8AjhYFAN0NLi9LHsY3WVzm2d5mYCSjljdFC
r9UwY7VfM/fZHf0QuVQ0R8EBbCp6IzS4vEq6nWh3kxitavc4MyedOi36nx/D2f1U
guG+cQh6098B80jtfdCE/iXccy8Rv0V0nRlAbJok0axuQSjfUQZxi6+q2Zomv1/H
GXzHbZVOpIdH0beouyG76ENArQPgnQ/NKwtXCIx+FVPifubzdy/sXR/PhjUmbLK7
Ty7WpyV5VyM8qGG1xAjshZMOHNMQdNiB+TMjMxaZjCnW62AjyxgC/mtGOVD5bdaW
fcMUyeoJqgV6rNaao4qjkAYtqnxNPPzKAipff985lZRsJ0VD6LdhskCNhUdTSb0J
kperTLJlfC0LNyO+OMfsOykOw4yVwf5VFONqKuDFcemXMDRCsO1Rkc/YZGjKbFe3
ocorHqUQGPCh84lLbsKg2QZ1dDORRL3PXc318agxZwyKfyGxCzMxZdlqGxAarQxM
bUsuDiaYku+7SyHnQ3c+OSvXAQfFGjTkUvK4J8qDO1B4TAeB+7C3f4XgfFs3lcHM
UlTRJCC+c3bQPWtkAeImcGFy78WW2+g9lPT+OezxuTcWWY9twVYpxACZ/EOI+CSJ
WbBQAYbZBGP0Cr2DxO/0QX/1FwHgIT+pGI7zmy7HwOJVnrC6gScVDliTsFdxgPlk
Y2O/0gf7jCR0x0iSc+IeXiegOCwEomTnm/oBIk+70+KXn99lVWs8pTRe+l6zoHPs
zCy0XLnJiodRJ0uicBIdqqhHiCBdSaHlxXJW10NRVhzTGRqxDOELVhHc4vGtToVP
eXcyQGAwTmHcogKFj+tmciQLOoR5M7h4V1fBV8aNk6PbmKhS9Y8MqRi/s8qRxKAF
22SwUIMMe6NGv4xVDquF7Gn1LK90fVhFtrDOdLWwmHhGLjBdDHYWmqHySfJCsJ75
tKvDPhML18dELzEZERDxh7ZrGG6DJPIZugKZVAW5FPEFYW7jozDMpH6DobVeBihm
Pl4DBZxeDZ+ZAbfocEm9vZKFJkyIDqf6aBSAD5wANEFEUGPGdEI8i4Q/OXKwG7os
l3mrd4fv6xskzZ0A0odwvo+b/GTu72qxWd488o6jmExxkQq2II1d5hQygDUuUxBj
l+xEuShkplsPVpDGfob1sK+Rq1zQEA3gBrfiCtK1F2F0HjsWjn3dQM0ActIKfP/0
8AzCLJumkhpAe68evkp619UB8HxLu5XMstnutMHC7sSfngHr/Rv0HnhMg4K9AAht
R6UH7G5nnC0w+T+iYGEfxlTx9EJGhGGe/2sm9FeV1DoTKZxaZuO7SRRswqBo0XLH
r712g8Kx5LuVZbeLUgvOZAtcUiVU8ZHDbqhOR0kNnPMOssnwBCTbmCwvJncrcyg4
TE4RwBPmpkPj11ZO3eoowKVFAccsNoF+oRTzWnPROo7LPpm3ldJLK7xP8liPfKJd
FT32WPpW68d+XLTYdxAu0ySFVMaE95ttPyLiJEME9PuZ6fbMifQebfzzmmkfSdvL
v/sM3B0aqBtYLbrtnfxk7feMfSPeLjQPZosWP9vGaVwINwDGYt9siGmu2zx2VnBH
cbm/dDz6s+SMQ4rynoBdAjSbskWdUuGhQDpNZGlRnlBgPKHAjNdGmpvL5x5fd7ez
3uAQXx/6LbkLH0ZwJToBumPgyy2tbMpOndFlJycfpqN81Ftgsxda9r1/+3tG3gAv
VJyOlnThc5Ehaav86q2yaporRAp1nIRwHicM15rjiDi303+nJ2Z28Piw0cX/0WpF
HBo2xOSIKlOwSzv4xlIfNPFBbsJ6PDOmWjAEj5iqZP8jHC1DmO4ueii0wCj9AQeb
xCIpQWppgmTaSLmNBIDdNU1u3y3PCXmKfIR/Vo40KZAFzGdzw9eflB0BPcYG89rq
GT9wzlOgXpJCoByOmUiGuN+KMcOtvrQQskxOMXyIBNcA9bBuVQjD2CQ+9TZrqqHt
bXKX25XE6idCJ+OmYK/GBWXHl9YMbNk3uS0qv5Oa6EOgj0Xz8a9mHKQPWpiGq0jp
Ri8J595fZJFtTxLKr1G2roTobYe+tYpz7CQ3PL4bvQ+nJGzKs6cMkFD7jgh1e5fm
3Af6t/RV+UAYGQVcfLwN40LDAxAokCsQWFELhuWmencykQO0o9ypLxYczP7To/SK
8B4GrW18a4mu81Wk7mk03/khC8aEgvyj4nzEQ4ALbf8/uuHmbTwKd+yk2I78mqQb
JUKQ0c4p5FEinTuYU/ixyrAr3hRRYx+WptSYYnB/Ha0EwDNwQovZm+SdXi7+0XAD
6tc/z39Atsht7wGc1YYkZjW/F5/0T4Zjs4H53pYo6xm6mwjiVlleWfdW5FAIoAEz
hZKVpLXf1cjxLoHq+TslM0oanxrpl9LofR9CgcIk/0feF0IbOw1OzbGky5kYF0kn
jDZdTLqHt1h9LO+am/fFi6nEKn0rwDDWF3sUdmubgWsMzbSSKzRIFaft+GKmk6oI
IHhkw49rsXYVgqb4b/4P5pavUJSENDbv486GuHNtXhu+BkAJxnVsduax2nQmwer6
dRIYr9a/J3+9ZGR9v15Zg9zMt20GATaKtYMyVuVN+p42GKHggbPwgMrRZpWCEgx6
c/BXVBpMzo6RpLre1n9J3BohAMeXmT1e9LORnsRrF36tRbcCimdPVv0raAnTUVN2
kgQzh0kB+Wr/TvtXAz1M/MGKXMgT4sGGV9FFER5Q42vZz9JHGr/rfvc86cvZZl60
wuWbpissz2oQr1TN3iBEWmPnTfw2W2EhFPxoTCFp97Ue49pKc0sP7tVLbDqhQ1mm
iAXb5bsxWRvug6nWYfF1MZUulPjHfhBu/2suIgN4MkKSLvGpjjjN3ptCJCGBbNIW
fiuK05GV2/kQXe3dGiFImtteSzE+wYhAraHa/npQGpxVJ4i2FraCuIhizxaLGM72
yx9vrgwa2503KYSJf0iz5Qg2SpU++hslvtZow8L1OA8FpTjqSm1qW/4LCakedViG
a/8b+T0wCcafSQFf252QrnRvaJKx7YAm4btbO1/kM+A0wICdH6m1HT3q4sgGimeK
77rPxeeftPh5P0LV80KZJIww94TWxoZOWU4iKN5f7GtzjNUxsXIwY9ib9YoBRlTJ
F/mbit1FscjATUQZwB09sjA1eBbDhWazz2XPg7jnOfssPSFxMSz9XDZ3+3U5KIrJ
fXUCWGbSBHvg+jY8budbTG5uNcsxPpnmSCiBLcCqXjU6DWjQV3ifR5sw7tCROPo4
WbtrHaKmzoqJObkyvIryEqboAtarCRI6NaDNqSxXyLWIFpPDyArmDaLezhk3VbOi
BHP8EnP5CLXQdSSP409Bv28pCtM8Ptd5qm1P6IsVI1N4k2i9Z3Qge9aVHUXBdjny
yMy5FjCIUJZoC85qcLHMMURtxJNY2pbe7FI415ugbPOk7Tk8wAIjD9mpJHFcmToR
7oopv2nqpRQ1brKGWaGiACF4is7A2xveJ78lelQ7keeGM3AbBSradPZiluYmHDY1
uTJBGbHeAObsyrjTwFE5xxAzVTpmv5Rq+pPuCsU3UBiAGuyZcmOkpt4g/du88REY
G4MnRLifOYt4OydOCyq9co0iGcFivzIaXcMwheLLSkhDZxzaSSrgJ9gp3p0JNhME
67CuSeo4tu6IZ8Bq83r6iyIfYHIEDzWXrSqpxRhtqUEwLaauBAuQ7z8lNeQptWpz
YFQ/wW6qqlql90ho8hHNB4sUcGxhdbZLqvVB11B15uAbYaM+Z42/WBQeCh1Q2mHw
b5YvfEHomkJCfsgEHcHjzADgWd+9q0QXAfoaVMqnt+2356TM/A19KQF2GTAjlQ45
yfh8RoenxEPWJXmWAlH8TLgtaH9uFwAMlyR0PUspsxaERS7OXs0OlKMLCQ6snE5U
nIwdrBaphS2W/cVz4FGejJQtk8QM88h/7T2OetFcI+a1IjRKw9b6vYtCr5CQx4zU
I4RGKL5MyEFiGquMQpoRZETg/d2wYeMrf4PUFQ2o4Ev5gsoI9hDTMOGGRdfjRWBq
Sn8xTDKIqhahxpmwrecxRH6fS/4WKFEosNuhYr9eN3USS6auvMZAf6X9TmcEXLu2
Pb6sNePU1OjvvUL9ES1Y8nQJ2syH4iziAChsBWLqAYZu32y8B3+zV0LNsTMOxLXz
GcZmfNm5vaFfwtTeCiAnKokYkPdA8bpVci0ZQ96+arY6+Co3jwRGrJjYtB+ZE9qW
W8soxIVKERgVWz1bcWKDiHkd7EAGwrkkpUHILZsZ/nZJs+/rroTtnheRDN6SabGK
rBrFvCzFbz+f5mbc+d2y1iVlLSmXIts8pcPhtqk1UxxG0LGsNL/FA1mJsJ4Pg2QI
1A1Q5gNRSL7Cgs52hxmJI0nY88d3NZTjMvk3K9zhK3D13Nqgw2bFNmeJQBJPJOKA
MsdH4saXRV0ASAQnGBJTh/J4tjtd2kKri2o6fxDxHjXGQ+dfY2aM1cQnYA+TYTmf
8MvSQclQKj40OCf9SDEkO2eBkmB/9zWWWphIoGaLJQ68Es47Yx5hgugahiNEhrBX
heiYLGE4NO2/o1DEJABPblINfy99AnrGQ8GV0HA7ZCSmZkPVpqYRNmUEgRZPqyzk
rivVnYdX/v1FxQ/x1oicjKj5pLT0hiymRJAFpKIKjkfmGxvHFX5c5c3ZzvZWsuiQ
lpz5NaG4QzOTvMbqrChbVBMixUVJba9TXmw/Fb1BcZpa5WlYH2hGUdyHpFFqHXQE
aOzpyRyI5DOmZKQay0uYaQnqqVvALrnYaxmj4EbFhbROv9ullAlmSnDALDHaa6T3
T4CLsHiUJMpwi5FtiEv/YuY3oOdbZLMJiXIHLo/VN3BLw/ttEiuL+jifTts0DQ+d
p5Jk2rwJkDUbf/8a7W2LdKdltpejZ6tqRqzcIPJ5m7ft556Gga56AGTBEjO3Q/ua
Mu1FTlXDT/EwCHvyZjQpjIeGkF90fh/Wc+hwUyBcFhfsAB6I/CglnciFv5Sg6/V/
izSHfCJv8goj0NogCFiY5WGd/Y2RHsrJJ8j8wC9bIKesaqHsfKvDmrQHQ0RPRPvT
XcVsyjiFH1ljjwYjjx7psjKsN8ugb2F8HzIWYV44fQWN/c24VXdQQDiU3StYXgSU
XofdSfyYTs3tRTgaoIuL4TRd2VoEgmWkj8YZs1RvpodqTVzG/SFI0n4uvEfqVVgZ
PSbxYTaYMkwr3yPeGbIsOkgA7qMA8b/fj9PTnhSXYu1LG21NY17dV/OXa0Rx6hjR
y8Inpt+EVC8UHbStnQDVgjnDUeVx4UoLy1PkV798LJSwEa81OTSPREsBl5JYw5nG
W4zY/HOqs5qza3TwjOHrH0RfQcNWiJ83eTSvI+7q3iYmlqX76t87L2o+w71OqiFg
/mlXRCIsYEsXuLyjBGslPGU2Nhor3iX+HShgsTRAzb78a94rrotiVU8U/VzVPfVR
ISYPIdNudoJVK+sEXb6/8RjsWa3oucK1FwM4me8QK8NGL7GqorRmBEf08NF4b3Dx
62h6czTYwWHB8tJioupO10+gqHE+mYju+WolI7Eof18uh5exNw+0U/KpOc90gQel
Ehcb+n7l5P+9PvZqzvURsrxn25hq8N1TGHsDhuHL2reuUIob6fMk8KcZ3Hv8lCHP
A3/vJfhz6hj8EyeU/gCepfL+EBe9sWUme5S25q9IFG4uZ4Rv0g4LtJ7591VdVvZo
5WsvI68zjzMqNpOpum1zyViEAD5+WvB1RE81xAFuUg94zLb4dJ8kKRnHhxbUwn6w
BT563IhOE+jhHY9ONbQyjgERV5mh3ZuwtLTdPnEbO0rboY7NWQGb4CfjdQp1FUBT
h8dWTZREIVgwOIn0+xxsLdWGQCFPa3gJ4pUeqd6yDTcdQQukmfGIiMZF4gv6rMS8
Fko5Go0g/1jxaF+aoX1V7WWR+bm3kcYeninW7Ed/lrrzDSo6fCPF6zrU2KdX5vuW
ZVTU8eUSFW9yM7HChN+/oivz5usQLYU2I6KOM3DnETSj+hVJKfllkiBoVOldnjz4
8Y7t4SUlBHF0LZC13M5MShz3NIfP4USV+bsGOV4+18kWwuSJjfIkueSOKobvV1w6
4FEIhL4cE7rEWwwD2i7xazyX6CILj274095hvkLDWEs46DSnfKk1z+dwFtz+8716
Lg2Dmo1kvrUF3uinKTao0er82wNIaW4PesB2yeZEZkAG7M8ng1Z58A5MOCGLZ3iJ
O4IcMp19GLvsJcJpXJxpoKRdjBoS+dFGAUAe4j+NdJLZafa3l/DHcCj1V0xAvL3/
B65fM3VCpq3NzbGEtJDA1p4a1MQHyewOe+RmOskzmGbgZ4M7PlFLtq36NGzY1yIh
uvD2rICTJF0ui5bBvpfBzoqaRa+OZ9AVm7zklXN06GE5WMVWHsdPqKSeIIqgLzm0
QGZ7BMbOAwg2Pps7fttyIoVsie28d3ZPDuSe2e/vJyEqhbE8Cudh9jgHPnXzreNU
9V660Gp4tsJxTB4OT1ZT2kWFb+Qk0tEx48QAUvY6GYkV6/Bg+AffpBPN43E2LvF4
pfCG694F6IvRfcKNIELbQlnSTfw51XCe6NJDDcjX1BBeIqzacXGmW+yMmZ58MyHf
VgQ3rWF5hg6Xlm5abGVjf33Cau9objoLBbaYb694305d3TiWcCSyzlfnhORMQcCc
WO1/V5ThnN2n/W3rgtc20cUpeZLNrgH9Qqcyl0cR7ZvcRsn1Z2DqIhbouW6s87hF
k+ujlqHX/7WjDhOWHlAXczLiszRdGoGJZBhR8GQ3WE/5KiDCbOrsvaEZ7uYwmQo4
yk5ZCcpk+xgMUzWg68MZtm3WL6m5wY/QHD9xSdAFBF5He3IR11va/3wg8pClU5yg
sy0WvQxq+BvOOr9QDkOCbpMG/X3MEkkWVntb+0SicIBZILbFkG/xS5MzI4aCXtp9
HcxrkJLkm8LWsGWXapj1v3zJrjR6ChqEsghK6Wf7wG6V9K6z3IkKyy1Op0KgAZjk
J+av6I8bGeCA6DSPlZKEWXGL/f3yC69NXotrv7MorBc8GPH1Ll/coEYAezRG9lMJ
gVfKM/Y+qppA9+cIzQP38Rnn57JrcFeWGHjhLPSZMGQoiDfZZTpeVhILv3zPdADc
bBXt5uHvqLXK11wh77SRj+HUcEZzrU47jhGrwpcGSZjRQOogXvuOfwLb1rgKP2Hp
wpmYlwpJ+Dce9chNtls2CLa7VHzcafiR5qmaYVjP38FM0qOg4oDILvw2HhidX9I+
R2qKAyGv0zMORaYiP/r1cxoKBA19fQfjNOat2HgyrYJKs/bx2BlEM1k/0CHCstwQ
9h+116soaZ3K7CRyIBjOGQuQwUE18BiSrT4IJ8JqJKaL2g8IhKapYNTe9FMe7sc/
x9ylx2RmlZdjK0oFkWZ5zKk9tNbFp+MvMq/FDnKiMov6zvuFfogyYCAIYrRa0RJ6
GuzmWHO9CKD3OeZhGJSm6yg0ObREsqqPYeQasYd0B4M7ONlDR4VTrr0LqA04uTbm
gaBZs5N9ZGpl4sSyl/zWnMFXjPW68JYlFkIsI6OWJUQRvQK0yaHb4n4IwLJT6bu7
JCVD3GLpo0qQG3q0B5Cxq8+7vpOzJOa5bK+kUSkXT/um8SeHaj4mkxnOfOI4BHkW
MzPmejfcej3dqbkgK8yzW4aFO/itwubF9/TJBi89Du76lw3dGQb28dMWjeOV4p2P
vzGONiB32qal/o0uYEut4QcKFQhGZDRS0u47KIUil21/kKiY4y/72xzTq6Akm7kr
dSW/DXyyUJJGx6srnvAOVCfe6hG09EcwoVjumwNqnIzMAwYivO90+o4bv5UCd1L2
gMQnMXqMp/sGlMuSOXFy8atRA71h48h53e5KtSrYdT0YYGDFMzVInNs5ZzLCdBHR
MAdpVnVdqu/fzZAjVQo8lH+1JHA0Sjfcpk8A46IqKjRWPp5xT+Lm5oabDqsSCF8o
FzPCQHwpIgJOqDKjueFnq4JO1d0VIurj7nI4shTHpPW4T1+AKD0BLiuN/Mg3vVeA
5p9BNNix0RPeazSsoq8J7nsbPe2jZYXzflhoSME5WqlN73Nxo6WJ+Z5SsArWlCjV
4ys8IpJLP2N9wqxaI0xaLa1PkoQYFLk0x5CJFxI1RQbzQ0EteMW5CxeITh/cBJr9
eLTl5/qpnt5Om0OS+cWpe664Z/LrKkzxnd4Lqll3O/fKOVu7t0+9Jr1JnVA/CWLQ
sHfFl42HID/a+RhQOeVPMxWlE+A+CEkExj45Magr81U4lixu8e0QH01iMAlCbA5W
PzL6KWpI3giH4ZlRmtQQLc97vkkIKc66JhQrWBp6/K+lkyd+D0pXvO4Y5Zz3TlEn
aJ5b/D+zTaLmmy+0pttmHxqejKacRDBJJkpsdIBCHV1BA8J+ZjnY1zYLI8PwAntp
YSCj7ijMXJVjjFUrT/hWau4Vmp4HW37URVB/EqkkeP03Cpkt+WqDvhX0uuH20eD6
48H+0zIQGJ3kk47hjiRwsRpijdy1TpK5/fbcynpiQx7YU5UmJxmV8gLLVM1vVh4E
1/HHKP70tj+T25vub2QFZ15PpXcPUsizfTGEujhC6TaUKe+iFxkiKxEs9I6yr0s9
HfSamt2WaL7fD6+du8R1znymXLNXB34ZhZCFRENeBeBXjHR/n0A5N7rDWKyfZFMa
deMoGNRx0tci+tzqtNE+BY8DJlhMBkL5o1ZRA5/z4E+YbYoUruxws0tvBWCwnl/K
i5eI48Z85qN1HG2rnGn8+qBOrPci/BnA6wOWmVL7OWZUTr+SN5Ecw5nHaSuFl6lI
SsS/1+vgG8q7aRiCO04OJeZSjor4fKcVghEl8ba06/Spou0eNIl5NMlFcjf+PUl+
PyQ3K0WcOTrsms48sFStft4TXC9pi45xmopt0AK9LfPQ7N91vSGDIJt5nwS4UpiO
pcXCs5ZTSMkmGVNp6ZYIpJtT2IXKJyGKBbcol2Mbw/gWoWeDlFnYqmSmfLnPW15e
KKz6SIE9AWOy2+9hi3M5yCJRBi5CYlAha9cO5t7Pv6Ur2pPzjl1yODW3fSDU06dR
uHYz3sTBIUSOZX4t9TIsRiTDbDBjwX4hBO+2lMSaQKFS3dOdGFzkXiAuSclvWgnp
8bGC8p+UK8lPa+W0wRDBY+9rCTDArQTNAEbQW6NFhkvpuqAU3I0bt8swEijEHEGE
QDlxRHzlzGUA5r8rlZwL/lQNf2ltv+znV3Bdb9SavPa5dbupvYY4nEJLOX6JMU/I
urZX9IOPCZhzYt5TMZOIObH2nHYXl8GoN760lXlY+6FqaI8A0UfFcZRPI/nwF33F
uiT4hMM5aIhHdzkbulJP+pZUOwe81qSuj77olnOIuX/mCeevcAGYuzNT+eITQOx1
QdvtxMP6nHwBnTN8UlyGiGFPJWzVfvd0yaf5AA22vRU2C7iZN76bFCYMlEku7oRY
r1otbI0zLQA0GHVEMsm9xJEJkLb5EWVCt5gEubpqoF/opBnrF80MSV1+hHKuRmzG
7BU4M90G7WQd9b1tmSt14EuYL2KlwFGkH9IrnonaAuT9dJ+fNAYbSBUnPD/lhAvN
iCc5sOqHGYO+QDStPwkd5n+C0yLG/AoAYVxxlBboZryWvfFhbUAumPXfdY54Y31i
BnwMR0ouP+e1ZwcMMqXbz0Ox0YOO+nCKJuO+50vjPeNGRNu3c4/8K9v2GSxrT5x2
JTgZ15EV7rYiadnpaHfF01CN2Nuyb7XQ9zLvIuAGiHEnSZxqWzN3cnb7RP9ESBVM
Fni0Kxn2C6AcbnbcgG1/SxkDT6O4LdnjxkaHssCjpV2Vvkz9qM07mGqHH8tgVUEa
OpeUURdg61BqMLKOvaeWrig8ZHP8NI6zuAHsE2ndMtB+XAQ2mNMCtCRq+YepGo7u
GhNAy3/C6Y8gnd5TuRgfT4qCIUtlk2TbVrfRqueDTKZyVzd5U6Na32IvT6YkSy84
3jIfji3tuRV1ieHljRbXZYQutKYDhvBOiI/yP8RSXO/ae3ciUDh7aqHa22etNlxc
rQVwy29+MxPTXjdY1uQ4omCgdorYi5LVGyysvEhrF2wqVDytcfiqRO9X3zBBE1JH
MKCtLm1Y2MQu06o5FvGMjOuhNT9Ep81c0PFTEorm1xE5aGxBMzVG0yP8QVeSOg+W
/Kidt5UeGjAcwJ5AEC3j10GZWGU1BNrL/J/MBe1a9PcvrugJmvGzW2CQWrskxuH3
CVK99T8oey5BeQfubF8VCcrsDsqOGIewyII2gqDSOSE8qLTUdoOCG1odKxgXrRHS
DYtYrB2crxTwUodGE9c9mPpPnXKGYDMIKcl/YrYlx/cf7nkCWVQPuCRHxt65x+ZC
LVItjGO9wR9RxXEZW8jxVXQQJQDan/Lw7iXAoZtqa1U0woqE3frHmT5RlfhKHZEX
qfsXLgvzCCvLNVpegGv4fim+pop9Ni3wtGeY5nrsBU3YAuhBkHqzNanJ9+n8wttF
s/91g2Y/feYaVEVsU9yJMaa9i7N5WtXHxWca854u346R121+T+4yVMw3C15gctMa
Kvnl1hk5tleE5uWY/Cviq1SgaBPxMOGHL/jQCO32YTs3adXqMt4L59Oyq+VOe17O
LFQ36scPIpG6zRPeQGliZTnaSgfO2Xy9CkeaDk4JAaSVRDfw4Lrn2RkqjQ79MRUl
JsN0hm/Xuivh2KXvmbDZ8Pa7UOf7O+VXOVTT6Vb4bw/pIhLJ0LsfM0MuL7XpRk1p
eQEZtMRbt3f8AUtaf5F7vKGMwoJ/B4f9+iYqgHtf/iR3rOXN1tL2QKR9kp4hcF43
CJDMm4ixmK4xyN/m1LvDhLB8KeWJWh9X8/WxInsKltUfTwcxUvpqVlrbf3QtNClO
f6O4rNAjzPLVQ6A3YqGbmu37Kc2pYXA+tbl88jehbL5Fk6wUxsDHMId39Sr+fQtW
e7iUYEcUuO7CtkIy0S11C51Em+/LqFtTYfFSorKSQTxIcdCHsxwd6w+4VNXi7829
YyXIvGeJ3mdR5njRMP9KiIZ3gCXC33iKOrNjMAo+AkfE6PRGgt+7woRmojoUUAsJ
nRMTPOPgdbwO6rBiP1UhBThdE73N/SdAJp3UphVhTppNLvYxMKBOArou4pDAuavB
kL+ncpFsifVGnRTzLZ8Sea7koxixhfrSvmtVzZXKlK3PygZmOncd9VYBDM4BeKqO
RKf5umN/+/nG8zzjL8VUcDpwROMZW0RpbRzB67GLk2XjTPTD/jkNsu1A9AS4OJgN
G9XP5N4So3pmYxxKuKoEKVhmkyJbXKoPO/OSowXgzucd/TJhGePcjk+5Q1jUFQ9Z
omjOcT6HpCXv4dthSgz4xMOsgBor19jnMRWRC/3fPaevyI00TWlcqDkSzABC3yRV
e3uwsbPGXErR5KWErYPG7nkPw964KHkUsUeJ5Mk9cZUZMQh1Awymiy2VkxaKuI/s
P0ZM2B9foHrGniFcMl/yLmsz/qJ5pjS9SybcooMhhhR2FPGpnkz7mb11eTppNqXD
Z3fBut/guSiCrTqpD+BJXSLq+eawlmxK+ECWRV1Pu7wMI7yqcDL9R2mU9AJTdPvO
so3NzR1bVqhlvt6sjD3aLjw6mdn8ZxMfhiXqqjo5nyAN2fkDa7rgHyCg/UdTEz2x
fKpmrjpyHHz85DoGfL6X4mF3pDRdPH4Lf2wRujlC8aD6stZJiHkVO1ZH2YCb5KDh
JkuouYcW4qNgC6SUTUmuGouGqbBTfrpaw0dJYqWIZsL3zBOP9bq/5feoggDAep7R
Fb/QVvOeRi11X2gAapdo3eIhW17wGT0pS8fGcb0E3fbt1yxLQWFKEvXcx4Fdm0LO
6A9GQKoSQDmy6piszKW8+YnBPLQYoPg1+BR/iI4EUJLm387Uv74RuGlcBuL4Aved
8Wtck5R6yhBcgAQaQCa/ZshgaoqaeYt4A8gevuC0HR/7lh1RuYz3hvmEmqBMIA/j
opX5dwiFMGNZCktlX/9HifTYdmnTcScTf/ZZOr6hGpt6LgQGPhm/gkPzXth9lJz3
lVPDZNqJGqCSTahHjnpuzujd9mWz9zbGROJUZ66Yhyl7KunWv27UaasvP5zzHwIr
LC7m946yZgrp7Cyf2gmYD8r4/GlfDST/ZkzzgFHa5oD99H7q3GM0fV38IbJzHOM2
jS9G2GWqmwnzjvt79VIn9gcHpZIloCdYVSaR1xeqT1AwP7RAX3nXrhXxgnc/X3xt
jvsMyTTF45o1HZ4llihnb9UDuQvhjFtTcJZR6YUW8scObbTvp6om7VKdxuKOHt/M
+cV9yHIva+CtZ6bhB3nXiePA/hamqEMjrQUXfjIllYjFDinrVaJs74wHzv6rQa2A
9Rkl3OsH24QfU0YAIELK+ULbJUWVnmkt6wMRT1qNY5QTriqX4YCMDmK/HTfuEd2K
er0OHpC4wTI7cQwwjaezHzfyHgDAG2MFqojq6t3LJ+9IU+ZHlFpOoH1X2iSR79ME
XJcEUsXPJ93ruErv2s8gIe45f/NNrIrGU3X3TVcQdlAIyxx5slhXogvYJ54m+kEc
IBJ0d2F3IBvPUYt3ZMUpA9B0766DJIFbkdlEh3nUmheUHX3DlQ4wBQcYYkTzcQXm
IyRNYplBxkeiFQEQBSWpbIPBYGYbo77F0wqL/OM7GHMsVsZn+JgcDMuLamHHwKC6
K/43048kyeb8NDYegUJZvtiOFvzE0LMWWfQwN861zDuGg0/zpoZ+IDHbDE8YMGRq
FTdCxNv6PJlGIE8+W20jKE+okJaNXI8rF+q5Ll/WMqvNo/ZjXXFBZUkgMCRCaTyB
smL1SnUAi05zCuC66+1v+DgtXb7Ufhf00HsvFk6ucBBTA0PvUa+n05/Emc8c3JAd
rXzoTyAa0ZN3ZdKnQsoy31kJTtZmJHRqotecSi6288AbY41q5+buwPSeoSwCPmB9
xKtVtvC/I9HrIENU8E99uFb/N6At+bAfGShgnvV3QuYtRBgNoCRbzd9gijSiio0Z
lswD4KAOuXIFJOimLB6T+up0DDNPony+DT/OyaJ2lsWLkcEtaSs6pSeeUrCG6gl2
0Va3CKg60Pa0DJg848+bsdPskgAEwyFKAf5FkQA4c88Lw8lyKKdlBSV3WN0RoAPD
zgLk9Tf/cbWNqByOWWCWA2wl9a2Yta4P9H5KEAXRLaQ91wT5hiAHKyWvzaiVZWM4
afkNTXMqFYjQKnk4vR9sSeJG6a/TimryEPbMG82pMZE955ZUoQ6Y2bOj4Qim7GoD
iNv5J/CgGM7ITzg6tBXAwUQwaOg8k78hXayB+j4s6XnJdCPWlUACIoGOkTRVDdn9
DCs0o6R/pXxqrET+AWHeS2/5nIVjrzYq5bOG6gfJBrmV0mHj0I8odq+qW+yWH7mZ
c6INvY20lRkji2DZoTtbAXFuAn1bIlmi0PZOg+UoLdVgSt/ieH83KeepqtGugze7
B4dryttPfzrGUNa4IfmxKR/gYLkl2t68vihefMvuQxX/KUQnpiLqReg2a7NBnYPR
YMdkwc2/R0z3NhJuHXh5NbRbUyBEPmksuYNV4EU5goG5cMGnj9hNf15/jkeX6ZEE
G4H3JCUJCnar8bWNNT3YRP4BWR2Z0stof38T0V87C7Bld+/90APiUl/7SUBX37Ov
Mn/osKb4BjBs+J8MGo/DwsJ9drV1HwUlb847+IW71vUgfB8caGqKvEoWd2kCc2pg
toayMA8tNZaEccvzAMHmAD0C3aFO8ZQHbQpUkH7sHWQNdjKb8G+Rjn3DoTEO8/uX
eaCyvaYrmo+yXtrdztiQQdDx2GdzjmUVkDwjvohCavGPXip/U0kvgAgUe/8aal5j
44DGE77vqe9G0OP3ezm3ZtYuXdTjU85Zxgkuyz5NsyKB7vLoOapyxcB2fYrBXdSk
i2ClOLf6YtV0vyws/090I6hxhUUy/g4JVgJdxEdP+OhVqv9Fo6D3BtSrIkA/WMQx
BygnYS20xWbQiOn7r/XKelNfgcV+aqVQ7dDRZ8BPC0W1+wGnI9tSasYwDOP/5upb
s5QxwcOxD80nPDflCAWY/IKzByBge41bFKodFqBw2a8q0fAmkjxLI4seFkLdcdKO
z8rNnd5e7azx6bMXf1s8BBrIjxIADA5O+FsZlXV14QvNh7x6todskmUou4BIDewb
ybXG9axk2Jaxp+lmNrgoqkr92QTcKEI0a1/H817ud8YkWBF8MhEnYfRut/H9hGBY
g014lOs+idD0khn+wmgtT00va5joRtVfuEBbRY/l86j6Kgqwtjq8IEhG1CRYPbCK
+r5TgBkgGn02fjpbFJsPiAo0Bd2yFyNT6/3NXpGU7MUWr2w7+op0G4XSlStU0bpt
cU0lT1xXpOqFgPmHDUr4Hp3yNLykkfmXFnTFQr0cMQFV20r3MrqcQJpI1tBg+sSM
mrufTC8zYagzWo5cQjeeEmi98eH70GkB9sxjektfCKJSqwtoO//dKqa6A66fTx79
agDmmn0l/P7sltOrT6JqC1zatL4wwChHbC7jMidtgEwiDUi2OdD3+GC3/ZuxJpgQ
vU6MGhxvbDkMfERd6ts4QFxuo9FEG35N8gy+JwCi+Z2W5MtKheAEgWYjcYhUkzOA
FJTol9hYfzbrFr3S965L+X2A3VS5/DtcqGqqm08Euyh+8f1TI1NOkbJnLhrS/NCP
0xpOKPc2eR0R2vKaNLdSPvUtPIqYKhizzdEJtAy66wbmeTfSXG52twkE1+RToFZ4
0wJjJSV4iwK8U/w0Cme0mV2x2d/l0d5/jwJXTGukYJgujkncdbplzAuPkJfm6eCz
4KnaUvgVBbTFpvpaEqF3J9RH6Z71oSTerqPrJRvMOFDNAktqdKz7lYOyypBg0dqW
i6FETNu2nVTC7GknDbN1xKmu861/nQlvslo7+ofwgmIIG8/pywtbYBck/W5/FA0a
50QHzHGxo+QftjfqrOMFxETEXrC7lNAmRwDb7oFX8PnFxRAmcVl9E/5Xp7ZDSjqN
PI408Tb9Wv/93yJVrWwpOdy0pM+z7tX7GmN4wpTAtwdWY9ImFC+hWBWEANnn8Ui3
lAGmyZgIoLDzGTnw+7B+vnDYYWsThJe8qTUShoSBxrZM/rpL35sIozOSQ3jDAWy3
2f1KNmMp9hdkVY8RgvZv/5Hvg2ijeJ/GR6Gx5K8fV12YmjJScJOALDW/bSoVr8gI
KTOOGRpFNOC7uMBHoFOE9MvvRqsL9AJErMKxUN8xsUnyfaDBRcDlSlJ/aXYADj5g
hfiVeUsATzb1tjiCmawlK4clOvCKMnBjetX10eUygjLgoz1pyX/IOTmM2SxKfJy9
yablV9lraXp6HEo5DndUfBo53+N7Vru5aSJuwvW2308yQr8EgfqJsT7gntbU8+I6
FwstE0L3/ECtCrovjDZCvgGEhq8zOuJ58vDNsOn1ZIN0C3qEGA6k64dhQpen5BEf
VXeRTwv8cKlNhsjq8rfu8Sj9atjUHxPwXyE6l+KenaE8YzgGGvygxbuLkgnxtQsk
oT86CR2uhohb5SobvGCwhKoxN/suYg/Wyzwl0JAehl3GjTRBV8Xk3qRIWUundTd5
P0DtB4ru7Hgc9e6aueLYMF/h1+9nktgRgKZ63yNI3dTuZLjnCs5geP6fz8nko393
tTIGDTOXtxBKX4w+P9sjUj+yL9nFn44COa69nU9qUGt1UgB6QMsEfgM8X55DbWib
LtOPDidJ9MttADcgDEghkRgN1hoRe7qmyp+syAbaALBz5j/K/tiid4Cp1+BZJW8x
yuzDGs2/6S+A28Jn21aNubiu9DR6mPDIkx3Jjlgk3cdu4XA7dnwTAjtU4vac20un
4k1eoGhKFDMXQdRr/EbxiyyUTzf6HoBBEP3nMebliRxow9Z8p62OZZFc3jAeBOJZ
FuZRoMQV9JjOHzXY+h9lf/wo2ZMqR+lUVPM4GxkKhH6FI+556do3G/8pkt0yAMpt
7RTZbAfF1Pakumqbj1g29fr/zwf793xa/gpJHbfyXa+ryN7ah/VS7E9oyp55jlHM
lL5hKqgYEjBYmW1OudNFZG8yiuj6Dtnd42knFwEA32qeM516xu8Oz8OyuulqqyRm
xreRehEeJYm2wNWpfEPRtEnQwcJ5HZn2LbSGodVdMK0CCV1L3R3h3DQSo4dDlPSh
z+oroKAAOo4bZ5rNoU/l5W8gtWmaakG4Z+AuE2iOU8BUH0U/7hXwoKhKb+RgIQ4v
dmptEE4NEYe63bAUO0QRUDCGbnwxWhlbb8LqMzG8CUTLIQn6GOhACoAXz0Os8qDN
iE50lidG8bxsKQl9FGrw1gtu6FtFouLDOSaFGqiTJeZfOLpv24tbWM6d6aCAcRpm
tcnssaHFeDvxs7qF1Cd0wG5Q9/Z7sC9mlvDL435dW+EFvAHNr5wa2AdNWDRdIaPN
29sh3+Ayenxk1JYaV4ag5Yw/P1Of8qE8QBVAXeLDXziG4+glgn1gJQCyPJogst1L
Ej+W8p7hVoZfzoIGP22UghP54MlT8YuazK6qyCvL8CVBSBLm7ZlI1W41VoIxfmMt
pssxyFEtUkpNAFW+O6WSLDOcxRGwZMHKWs5qw66PLMplzA9e/NGUbpyhEpdkZkUM
KtAVBdIucJW1BSVkiaO47PFKvl1ZHATDF/nHQENOvRQPo/EBqF8XHF2h3RNnaRb1
iBInFVN04oE7gPIubRdsMRP9ItWE2EGHUzm/axaCphZdJR4L+IA4gSQvf1nqvGgL
khUU26FsK/4R7hCmHUZep3aS4YPI/jbyKYL5NH5hPM25ytCQhH+G9756sa97g6YM
AE0HJR+juYSf2KOo1BzJuMncWD7sr28Ra425K7rLCzfSFE490VhkkYFrZkzFkF3h
qCqV7HwDZzBPpm/RhmjJI4LCsVk9DZobzfMmo+OiPGFhBFiFjXJ5GX5z/DTgJCV3
psNhr3w68bRU9yqb7WP61Gl68CYzx3GMzlSfqhkS1ImxsnX+rEpKlR+CGSkvZkGe
/GZnpYC+ByXv6KRdPAeSkbgpmT6ty4m5UctqshGKKejDuFozI0ljLbefY40wXsR6
v3VH33Pb+gX4kdShqI4HGXpHTSs7SL/fbpd0BPgduArN/dQ5DIImLURDVmWyVQVj
u+x8G2Mx7QsFlr2hh52zaV0txtaW/nlr2N4eNwQVOkdp8UJFZmt4gesEXBh5Vvuz
0PoQYfoXnF0WobsRza6C1sAA8BGQ7ewCFIvfEadeNF2IwjJ0ZVvuRg/smrUWjuSX
hfn/6ATgLi2vr5fVrw9OYjt/MmgjjiJovoKQFlAW1fDra0IEII3Cs2jaEUHRnj4R
tBfhKRaIAll1xIRerd2E5eFzAn94OLBbuCXwz13tW0tUqm1qnqBBF0mKrm8rhJsR
TZl0RWnfiXxtf7dNn9T0QKbR26Q0rTYoWCIVRdzVcTCjI8Sa7mJiFp6ABuTe9LUp
FnoPcEAukgjp3XWgm419eWlLkZ/bFFsgX+FxcMMaM1tNtOnJLPX7NyC364f9S0Qx
SDFXZ3O18LNkegEKS9AjNBOX65RAsBcKFGrT3QYO07Wol6ugpeQDLHOoxSco+tad
UmQ0W2/Q9kNTi/rmqHcFwNK9RrFfVEXgiRIkfvBvnIbuy6mUQf1RfiDf6S++xUol
/RPKAoKvATbMbq+y4QMNeF2oALIoKgE1uPTxB/4QzjgwhK2zWMCzFrhsYmxFPgEp
SKm5G/pZ+1f6oyTEijoTCDavnnMyAN4MjQ+QHHKjW4I81JPxZMvO1l5tv28sDYK4
ZzFC/rJ2P9hPC5IWUDjUsgpDPTn/J3ugPW/uSSoRYm9uKj5hsZuMqwz7HVgW5c5G
1Sc+UUzZ9F4DHpw0XGVKMFlwEEOVfFgcRkZyiXjh13MFbaDSymsJMF7q4nAG/jzL
xWLqq44pGPCmxvpvo7DzhsihkFecPwvUGDl3Zg2G4h2e3VKv8oelqpeZ8oL2iC+5
gnNPg4oe8irZ8CrvELKscfPYY+2BqEXx67uSC56zQ06TaQ6kAHD11vqLIrtO//37
Hbf51aejlv+Nth5GRj3vZ5omyYYvglltkPBdmKTbPT+NkMWyrt/vxRebR7ItPZQI
XitVqyGKOu1G7C2shadAHKNEbG9eJAB2JJ/H+i7TEXIReP39NYbk9/wdBHNabouZ
7vAXKlT+n7b0DpePSouTQwR03L5dbGuwIhusKzyLkluko4H1qf3hKwKFE/iXaOin
DjaZD2bVfVmIqi4hr+n51C25IsvMjHAzWVExVZB15Pi38pIBZAOtLGwTMKs8Sfo3
xDolbISIQQUFvaFoz5Ovxae6607OJcy173iLKMq+NVAF5l7frZ1Yu2Ny6tmAbg4S
LJu8IyDQnvHPhhiv2ji0KW7jSoX1+pws4QPofSqwuzKXpXRWDTMr1BNGWvqtrgsj
If/kMwC1Nxdm46jF//zTm6ATccwNMRxkrLtVBxRXt9GlWAfqSOiVmcCIpcTCJSOQ
x7tY7vUWhoxKwgh8h5SdSKxJ5wpHfEetfQ1Il5B64NghWf3m+oi6qTv7FvQbIK4R
mG3ZO4kafa88he22ZM7tROusVU8k6y8AWb5iMhtB9ENA12PzTI5WzdW2ekvGzb8U
VTnJftnCVWq5s7tuCl6Wj3T3XOHKv8L4KA9/CViwgQ2VCCMA4OgnVs1hXsMaxEBE
FxeKZgZM7OrymoKeOAzBwK8wLFeVOCkoDuSxAqKIZnu39URq4YFCcsEg/EBijWSi
UF3zMEL2WrsEFzgT5MARQzJxE/KxoJ8bHFxSvpxedxF3HtYwwBr4YQQ4Yx3NoOFV
VvBuWXVjtJah5MAc+ooggSKE7OK1xkJt3FP/V70WyrgDTVOrIIyFWxNvpeLLeVm+
w8fQc8+LRd71cQDoh2bkro62Ti16rd1nYa4n6srqh4JwsEf2EaM+WtE88Qj3xV4j
JK29560vCQTuB2hLzTc2WXMFzgSMglDYF3XUauJZzac04OPlZDOAP1pJDrc6Xznk
1CC3dSRMosPZ+Jp7yIgFd0pqfFQndMX+CJP47EkA1kkpMwKejnJQwBRiklVDrE26
vfbYESTaf08rAuaV1gXd6/CMLsrgGRhTDtVb/7JZByFV6GsAkBsNTehJdxU9DN3q
75R5tsPj59oZdLqnrzqZcBr3S2ectjjKyv0tjHsfVMJPfES6/BJaxBnoIJZYqAqC
KvJqf2NqBupb24WUux50aik4JZujNuiE857yJZNNS1Hw7w8s13pj9zVPfv6jjk8R
CU9RTtsGF05H+u6On4lvuUseQIzGpoUexMWcXwwYZWTidQLZZaermGQ656/vhSld
ydOg/o3u/jdlsLFl+WX9XX3uK5vAgRvZqPDPbCqD4aVGhzq6KijF091qMOdRKI4X
KTFk8IxchrXUFZnW/SuAVbu9XCg+EsfcEpsQiDIYG7nFB38UPbm2Ri93FdFbOeI6
5hHU79wB5umfQqRUQDh+Jr0QzPXQb41Kqwr3CriXxWuTLYBKG4yR+H5kWoycwsm4
u64cQ38xvClFAVUG4x8PM0AeNtXPQSKmuVCgfYdf7VLQpK+o/OV5jN3yVIUPloPq
WArfj7Rdoap3CiOImT7P5Hz84O2pQ+9JMJ6rTzdBu85qN3He1YhvTEy1/SgK989s
M7XKCPWh8a3BngpdMxopbUaGo/E6aFQoE244v/tpWR2atpLt90bdLV8fxzFU2roM
EhzJMd6Oza02CyQZBZOYJ/TlXaJIYRpXdbMM8nd3/3NyExv3xeq6Z8wVgeqZTMS8
rFOXXdIrGX4+M2ctqKHXMyojhJJd/8e4oeR5OfxI2qUsWE3SR95XNAc2PlEv2Z+o
DijIpEE7PEuRECQ5iiU/8RVvlg1ZKVkEZDC6P8hOzQ+dEwvymipbWxjVVDpCaxQ5
P6rSzqfqj8M+x0QHV71d5VZpNUI57NCQ5JaSyv08HQ6PDukSQ5lyEasB9CP5VX6X
PpzdRFxX/uxj2QNKbHL17e1Jp9PMoWQvyOuOyy4wKBRFwnDBnQZnG/ZYPqz3jllg
4QWI+gGcBzyuNjmASAZfInQS5iL89tkpmKUYN9V3NCLSC+RA04slmUNzmRLGVFEb
COjZD3afLv2bFfrW0VYVUT7BtxT3rpOKQEFzC8YIxx0chP50yMq4hsftJt5Cslwf
gEf4pBsu8A+1C+4hqFdnTmUqkuA9L+hFVpdOl2udG/xV2p2qGe0vCtXVgOyJhOgm
2+7MOhvc2zcibPLh8AaxQeHLTA0jEL5MBa/zzfOSEjkirz92mjmfIRjSI8+VVK2F
A9g6G5pIhQMxhUBg/OhFl8fXLrdtITzALptAy+v8qJBa+YaYxs6wOfl8SI5xzjUI
mCcEgV3BvPuGuNcsN1eraOyou3DYx0v2dGecT5XuBJRvWgm0d7a4gdVbBWDCWzeB
FD5IpKrBit75cEBENm9WMpTAJ+iea7yptsYaH88zPGZmM7kZ8jXEiXK1cqa6+KaP
/A3JiJ8TjaMyj172WHCrlcqiDZSas9l8QrMEa8wL9vEvUixS7O63eOBHSbkqpVNL
xTRmopq7wACHQ55E+80v8rQY3JswkYh80Zr3Nb7+fB/l0ArBD7GjfJKHimsgCL48
s+RDp+ojysTxsW190m/Y1lfY8r0zYUqCSw5oL8qiutxPJuwyTAKrPVn9RuBMj98O
zDWKT1wEP5Niszu3eagkP612Ym4oNleH3eabpe3M5LkZPyKWx+QCpWljxXDBAib/
HixtlQsQPhakNzWG1495E9naYpfnLJAFMDiHGZyrQrieXP/87LOXKI4G2A7rcYW6
mrLqrrdfQ6KNA1tfxt/wwMoUkYA1ygS8kVOJY0W2V9i4X0ahKgqRsiOr6LSHSu5t
T4ciAsWRF5Zhp3rjPcxIxRT7KqaZD4gnGdlpwZTTA4+Pk27+4PW8CCCEkYUyhClX
1I2mpZPXOfwQ0CvTEbOiiMRBiWLoR3upU2/7BBzFq+xw/G974Yaf+lumaZzk1O+L
fmFvLoQwA4XF28RwVqSB03wk1k7njmLWf8SHY0Psnzznj/+D5IP+NiUDD5QlyuCz
qZXbq7zebGj0BzjRPmKIyOJJtdO34rAmlwIiouNhWbQnXgaMWjWolW6cnyXLRDFo
y/BKD0na8KgM0jmtvH7+1/j2Y0oh9G0Ctignmfvht3r2KpxGHbTVnSFl3tlyGpkV
Slc3KzGELHUtlbZmbnsitNH+7QP42wh7zI5kQbqkbJ7DxV8r9YY8WrMovjBxNiUi
yUgyLc06qLXMURr3YShn22K7XfdccCd3+NrXn81DGl+tziiwP3le7VCGsTBRagYD
7KeIh46C7Ck3yZasIVEHPbcyk/Dh3A0pytMCQfkjXqIwMoBvbSa0pYG8oDMZoQIW
Q4Nrn6Eik9V/qF1QJXmVNkmnRGRcMIcxIem+spgVAZ3JPWqjL85xKrW73sYZCmEa
sv3b4goFcd1Llrc/nCmUw26OA3/Cngj3JCVUwmq3j897wmzq+u8mPnVscb6vRUli
CDWMmkSobmrsTGScJeQdGc7z7Kmb3HjUmmJZCKJXfRHeu+Manofh/l3OSfq/8hBB
W2vYIt05HxqapwMRf3bw8/ja2miO30NmrHvL6+MXQe5PUjMO5P1WNOtX0i7CVVNB
07ym2hFUM/5yms753UTN7PBfebb1yW2//v/AvguWrSSNXBwxR3cgKnbAx2v3KEoj
osjzG+NkRei56LU9SpBe5V8d9QSzT+2oCGAZV49ByroEXOIHGW5hj4LDHbH8RVvE
JNruRc9X8O9BlRgN2ZbtYy/cweKkJq80doBfXPHWTiK6Z+YhUeTsNflb1sJivahV
IvbxkFYCEEz2htAQIsGRxFYJF1zXpeXltK2Fn3WX3Um/Bk76b8s8cDgEumHy4Stq
7O8PPKlGtAsK/TKUeh1967ygSuqYe5BYfHmYAT2VwxRg/llbZFQqfCQWr0wPG3hi
RlpqPQIE4OrfLD26nRtSjNzr7PhYLxW3S0cFcQ2fX047syGYpUj+5fTVOUBqfbbH
n3svNc0NwXFRbmSKuT5PeCgCs0sAzjKpR432IrP5UJjb9N7/7Nbk9sHsGcWzKiOP
24z4jIWZddHKn/olPBYt3IEhnTxQGW+f+iFbR19nBh+thktaPMnCwZHZs/B9mE6S
bq3I4RdL49pXhDFE0E2vYS/5F+DiNH9TF3hYLeyA7qVxa6HRWUcZHc57EQMqwwgg
r1L8K68K9glLv4a9Zs3Ui4PEDECGF76e/yzgWwa12IK5YwR7PJ3AXaYPQ9T8lAYm
iglOknQ0Lmqzfa1KuoECQ4VR30IHnCb4Rk3mQSC1jWOytpyM+dglfnjDaQ6J++S+
fTWh9q2f5kAg35t5UVejQFWGUKWldZlNdb6ecsJn9iQbqYk+7NRcead7Y+VirbBG
S0CJPDUxJ5DOHkT5raodIJL2WeEcTplomBrPMv/rrYf6rpAyn+OHHNPylxQjhIh4
moijVp0Fs52svYvmd9XhHUHIwDO93Fayk/y9KUqlGr7L/Mf20OQBLZE9S8CAa7hZ
ReAwOcv8mv4HaWOW60eAcr2VxmYPiu5geO4SCjLYc5mye0BC/7cGoIi5qgagd8pn
aYRUiZjgkDZ46lEs8CP74mikeCzvFLB+3hhJqPetotNUF90/JBCcAnbWvNT0gFqr
e8SrQduEza4kVx5oK1h4u+BRfBJaikUeVuIwZk13F8UAslwkRSzO3gdWN95+DQsr
YwtviTGuw8qXVY2f3gAgqbONKlOBGUoi/TjthB/MWZA0Ijbv1ncd7WL9N80Hc0s8
zg+Psk6QMZ825Kt8DC+nHpT889x0BC/jfyqi4jqBr6eCJye0O558jzZTA0/HolRx
/NOoipl0IGdKdm5o920tSz3fK0mk++LoAaGv602quC83poeDe2dMf/lGGi6qUjbE
1u8zukk6OSRL5fVMkXYfh8yhZ0/say8cITg74dUHdGsDFoBlZPUbJwAWSWsykHW3
/NG3bqar+qIii4q7l7hYqRclEOYS0Vu8D26LE9+p6EAVEKZROf5UORrtOgYqQqO2
imhmUTILknEKMvPYZhB/aqynadTjYGwRYxbHLF3sAHS2p6HX4iNQSkPKKoKJ2HsY
9wnMTnuYeopyPbZGggGp2tLUSGPVQDD/I408e603wE772VIb39dNCmBCSmezWVCG
3ETzP9aXR/i5xhZQwDyPptXnD4+sipQ0UBoJAXHTzWihyWSFDHZQunTVw08PB674
6niH/RNelX0iWkvCsoc0ayp54JfJAcTsykD1eChnVb22ZG69ZE4LF/6P8MBiJxnk
+5qSbN/ljcNkUr+L0rkFhfuaS8ApowoHvGdDW+s2X6NSLbBTa0rfqr7bzb4LR8yU
L6BbMkU2FbztuQ5G3yTMp3nAklsn7qljX38KjUVMVq4JbeSS/avSa4b8C6GDxKkH
N1Cz5WQJeHHFgpRSXE+Eh90Vb2pEMnKlC7jey6Z9txqNlyuLXN+YP7yYzao3Yop4
FldzPxuPUd2xhOAJPvijfHpPOrviRIe68rLXjz/pEHZx3q9mL8uvvMNXN6d32op/
mOT31LaiyD6ZQxuiPW3sTAMpuu5xp5YDgP2fVYvjOfQ1SiYDzhNko9bx0FvfZMhq
u8E+x0NSN6XzNUe6c5KJ4BVC+j/1HTGNfCsYkunnleGZynG51K5sBgy6+q0uMbFo
3V+Pu2G8EBJpZkS5OsAV64Y0kDHRZ8XrytKVBxoAtNwquKBeBj5+XO3FWtxqEF5G
uXO5AF+YVbaQYFEdvNF3uGUiFfHbVVm2bzch5ZoHLPKymCuvU9BKe+lmdZXdL/kO
22DfsoOkNAIRR+ORj92a6SIU29av+IeoNJfui+COtA0vUIPStT6EB8nol8CS3Jxn
eIvbisMi1nW1mu+BHBwE1gBCCXZ/AjSdZvIrIQRMegAcW0etRvn+qKG4ajilKHWO
3mb0wWEPpu7e2wjhmxUbOTSZR1He3Chpk+t3kP7Hhq8Fzhf5o0T1UUkMAIn36IdN
YVfFMVG9EIFDwMrYHOpEyoCo2OuI26oCTTRo3PCnt4Bnwt9nLV78cXNgViMKcIWl
LjN2K7IHyooKR5UuHrKq7H1WzeysZnQH/3LCfMsRXUOFXhZ+6fWIIneRLiFp9KAK
xVDeDWTTpBAVpAO160M3tI+vskI0hj6Pt0xgkBWt+kwEnPHr2RNgMcQynTr3owpK
N+2yMKmsthJaPCwujewCGyUlpUMGGM4NIzGLzOzVijE0iQJZhg2K3MNTqBLxcWXn
kGlofEwY2dvymABkSamtvVZ9gqguhRhl8os0KolfI3utDuHDh9+HN5uzE5eoNSCe
PwtT2hANgPvCnBuoTFBAI5NyE5uQDP8c5aCi4aZSZUXnYOHY7wa14+tSvW1AnNE6
kdMo9J1qevhf3pAGOU3ldElsGWBh078Lnrmbx7/1ZajMNuxBRc4zSvoGhEhosKvY
zLI1drbtkWVPo54zrdCL+LPQg61uIOe7owr1Cv3zFN7Ja11Qhil0f0SUb6i5OtP9
PVV+1XxRXjsvwHEGa3LHKzF+xY+eAX7NtxsRKDZza+WqurC6CaYF9Ukapuww9mKC
jtWPww3Qrogyd3joLTE49iW90WJWhs7y8NYvRbFn8RiXSMyRdc6HlxpO7/kiMA8H
gvNUyQOe9dLm4R93OtOIEecqelqw3sA29qRfkeWbHY0VbDARpJ5NclzmWBiGCZkV
9UJKwFVMDuodFTjpsQ6tSzuRvKn/8znr/brl612eXvLLOeVoB/KbBiAJmEecS+9c
M9ZcJF3JLR0Z/cSEJAohibVRXeyY2lPZzFkyD8tVa7Qx9qSPRNBUG6Gk1NUrY2BA
+1L1yy/yN6isXCq2hkpuBTth9PHwICruNVZSFWM1o49HaWxnTaOafHI/NviZR3VJ
+pnFB/dH8SpT/5eWS/viLVHiXq9+vvPGNNMOhwy3E+4r6sElby2EqtBE0ixEiF/a
bdYxY1p1hwidFR1wI091XBfmc80oVzH9eMyhAYroAxul7xTUee4PK+EVufVKdMkM
Su2jbPzXz11gjjP7Wte17McB4G9ZGRJ7i32IGSQtFgF46Mr1JqoPRQEXzrpA/oc/
PrcxPGVEIevxuckGC7IgmkIOEpJQJRGvDJodVXy1XCxLkGxGBcp/ioc2Xaqnr8t8
IjnlCcREUeqmi3KVpFGPUkn0PvwtM1eaDcQJgrelJTcjJAzoOdMu9WCRcTVm0Yjt
n+Pv4db26TE9b7uodGIJZObT0R3fwDUBs9VCAW6/2hAQGcKWDYIYmdVZZ6p2uyyb
x/esW3PyW+7XeMTVZyJBoCF+TWgB61qSgLCsanyWm39v5kGG81PhHr81rAOM/xlB
8MALi+hDMfTQGztBlLesl8ufW5gkEXrOGODDwyDwausy7mT/PcdI//72Hh7J22Rm
FeL3lrXvVn8SbMODy2tRvuKmVQ7ny1Kp5t3umJq/Bo8OXCn+FXWnLrQVe+bf3p96
I2lz/csfCZBgo7UsifOTTXKFyf57siZrsVqSt89oDHGDghh/34D7RdbDIEytA6Fu
Z8LTHgByiOkdkxS1To3QteGayTVAGREzP1PmINOE7JZD9Tt/RJLvctMP2U7WNI4Y
+A7r52qiXo+XVT8zu+lkMb40ykB/6Ji1UtjjAdsGP4QzP5cfNnU488tWlyPO1Il/
oix3ALjXTzSdYanMjrsBnfsezIxhgMjie1DfNhyPrRQwlLRejDxU5DcHh3mEbdoG
nUIZougyQmbY22O8YGGY0MpntcpU7f8Bi8qEclfChJE+V/58EQOSoK46M3XWhGX3
FmysT8PFfWkhF94CGCl4yHOsOSFfGBfesuragEtVxR2uOpIVxxgieKziZ5w2Wx4B
MRGCFi1LobtX9WQH9kVRP3vBwUo2PN0Ed4ncluXakDlAw1rSKJ27LHaW+hUFrBuP
yCAPjcZxraSErUsfJIVYPLZf4H6YvcrjAlaOqMILyScbQ2LwtIFGdbPC2zMlIcVq
icDklhenHiPRvU46mJI0SJuzEBz7oJJveubDtp9Vf88WlSCB251BKvDlO8Lid9f6
pm/pV8UJs6Tueu9/mxGC3IXo1LjCdAIN4+IO/Y9j6RakaQI1bPoq3pffth7JUNRZ
/88rgEw8vAhdVGFVkH1oEXJb9VUiBdaqM0hqGm/YSkfzhuOykmU+BDF8V3NnSFRE
aScV6eVY9omBhXXP8O0f2qioJpC7c7R4DUoImbjdexNs35JZKnVCyv7+cDf7pXVo
nU6ENJ1gm7bwyL/VNk7rf4q07JygnS7pU06QZJiLAioDapOzHh7ZYPbJKzalcB4J
BrEfsF966pZeYB0WBwklwDwirEIneAYHrSx1CMq0mItljSXWIrLEpojh9iZ4eelG
bKa6d+Jm/+4l0GA7MqDpkAIi9P8y8rQdlMvk77plqekYZYBJF9YpKmXQIIF4G4Wj
y6AZTKgHLe3kpWfPaKlxpEWDnmbzfeIKh+FNsZUR9PE9ZBAlXnGBKiSyhIecT8Rf
2UY3upgNnko0uf52svOYaZYneqSEuescYOiUBOGo5XghLJi8EONkO7bxeJRXpjW2
9DIiEgOi09oHSrVz9m5Wx2lTFaW9b4IplQ8hJUlpzrTaiAkpIUZRTkGcnWaxlHO3
QB1Zv0FvrzQJGtHTmRse6DGNqI1z8zTF9bDfxTcX8Gm3Sk5EG9JRCbhW5gZK1Us7
YNr87ZU/JNM4/5QPXZML7wNG8nNQ7nRJmNlVwQ2L5Tnwj5c2MtalD/I06tibEfq/
O8JpNxsmQV4XMiX0ByIqgBQEdy1aYtDeEZcTrX2TLbstjahzZoZjbWEzmIX9Yodg
SxlfH6zeLApvvKhvLVlQUno9nYtNbHyMGfb92vq0PUwTNAAMkO79nwv9bWX4cWLo
nfhLWwQMdx5B/og4ZJbcSg7d8tOyWf/5PQSysR4ZU2B2Qq+zZD6lgdxzeQfND7do
LDJ648koqP2xVpMePLLJKV93QFYsR8+BprDJvaVetNZPQxKC8jMyCjs3AZ9LgXB4
sPSgyKRqzoioWVsMxg02GsQyC1QQ5qsfF4TKRMw/VF6aNGlUmmH8JGFSVHbNqWiD
xN2tOkMqAs4La2YhUbRYBtH2y8VlRC+NofF7lUSDIdQSDofwlslRPXLzm1TkXWhQ
WfumTtsTlkGiiO3owv0+LN6lAH/oSPj1JimtMFuKcqM/5k7M3UF4px6v7SaqX8vX
vcdy2ijy/wTP/jMkERTdCBOJh3r3bbyvmwJdrjLPbgnUp0a5+bgYMbzYYbbHRPqA
7tKXrISoBiE5MdPJtQNnPqcK+JXz7CarCt73eq9rGYVP3TkfJHTzUZD/aGZrlhJS
LdRekA9dOWO5Co3gnF4ZRO8iO75xB3T0O8odPULFuv5xsEMYFQb+lcDC+9iwmVRg
TEEQxlwwgFyhfR81AMcFTuZzjfjmdFchHAgZw0gUPbfJbXAi1dPyHGJMAcqZDBbZ
39/LeixMSJD+ReR81pTqsTgGRC+bqrJrsvDkS1nK01fdYvL7X95BdQpVjBu7HXsk
dSOgXcM4/B4TONkun6i07yTyccrx9w8yiAlW5yPOUCw3ptK1LF9erGXxb59fgxTs
SVQeSuP9IOPXJanfYDouTXwFWkjiUnBzrQ8QLdLTF3hsT9gt9cezpMoQoTO10P2d
3/QahzyUut0G2Uw9YDK2JsIEYVx9IgdyJXznAd+WMJtIPx9cACfRWnwcuG7hzelC
Jtuoho8d2j6v1dFW99AibvEyVGXW3yuhRhwQOaWhW7iaeqPZ6Twno6BhBEx4ah0D
IDEXSml4AROtKL1Sm8HQhdeIaXm4+W+tXQeo2Dp9T4JV6F2kd2P1jzJfN+oF2d4Z
ExDGDFniNSJgruvzZ0p3iSSrfWbTr+AXBXJKPu6WGAPDVYw9SZ9Y8L0i9N9ECLmu
IyHFi4ltmA2tQ2nXa5CSMH4frLglQ3hPJUGflwt3CLzRTaREJt/p+aE68CTkNdEP
nN6UDH6EUuN+CjsHFLENi/6g10c9TEyJdaR940Inv/UDEl/LW3+SzXDOIrAmAUrO
QC8t5P/kSnwcl50R6giDHU/cXvwrlVzj7FOXniICNDZ378zllgY1ilIRBq7MZL8u
G0dOBUfCbSd6o+LRtA8EDRCSa4tri8bRanAg7nj1r5SzrpDaCOvZk+5XASqb+Xxd
QgdXhYsmrDYdpzGXNPPPKcpkzkrQKonw1wvrrimY5pJkNhZMyEVA2t/ug/k2BDHN
AC07zvmDZZGBB9I5vkhVdSDYscDnhjuK3+rqrUjjqEacgoTEZci7Y/5rTc0Zr4MW
+HuyReIS5Gas3xs9vVGVtyspBydLkGaFhf1iCiWiDPeT0UEsKnkBBV0p+iy1Z+vC
f58h5SNCBTQLeB5Ax72JZ1k7yUYjfSnSgvnMm1XDoyD/7tcVRXdOT/VhOOuceK3q
F3JNG0y+cj46ZUTgqhvaRTI37QwYWhS9NXInaPujdA6aT1qvHi0vU+XMEO+LsKFK
eayNQiswDSpv1hMikgKb8YBLDFgqt2jR1+xF+XuHqNoMi+Q3EX134TdOUye+cOUY
Ui4ajRhPj6UZJgwVu3+E9oXLd5GQcUdQJT3bIfiEh6zCZKQBCk/Ih9ET3rnnh3/w
wjtcnwpamtZAOopzNMpW2zFfwQbYw7/nLr0kQA02sq2q8LTaXWmXQK0fJRNkbiG/
dCQVdmefvwkjc9of2Eqc4TWSRSj61Sr1c2Va37ranKgXnO2Rvkc95pnQYto6lFKg
rm9jaRdc5OtpCzwHZY9EjC0ZR32ruPQ3TlA6sD3SPKaPYRHthXCzUUmSkiA7lwKQ
9HndZcU9zI9hc5OfCXcghDMbwr5p3ZbuqAzGnnijuWvqnJnbELDdyDZXSdBLpHeU
NwaY/BDBoiXo4e5EaumKmU/fZbquh+VBX9Km0uX0G1UrnmeHIinwW+VOae+Z0PTp
iUY7X7IJ6/34xFVroO9IbavWpWeSLWNGJAY0lojACrOKtjgoqlZiwy27neg4NCzr
Xm6q7TuWzMd4CIKwPTp2n1v7LjFsS5CsH3bybgT+Ru72XeEUW8YtsyBGCnYM8BlQ
cMZ+enH/fgONEuoSijyE/PGQq9k08NTYuFRdvfmjw8BkhYj6mcSNnjYRZsB8i75/
hRSWdEFdxz2xYgYee+nR/Mlnf+yZc8hxc6vl0Dc7ryvMJdKjNyAM+Pa5FtFZcJmj
MPmnNpD5eAVaE+gGG89l//jTbbMO9DrAW1eQfwypk6uEvCpZB+4L11vV7f1n/vhd
u9Si86u8nxtUgtM/MFTqx3XGxSjXlWh+94rbgpo5EKN+tIWovPEmhf/6WsHziknW
M1KGG6VI8fj4m+l3/ildHfizHBXrLnD4aGPKptdc+CusHVslg7L35P0b7ZuWygPp
kXpERmFN1oq4QikITvGhtV6PljsHxszyymRREzz5vg+vswGuFE18Gf1NVLDG431N
IhM/u260rfbeCmAUeAv3g1ZXjLt/+mQATgslEdOxiAzAFZmzT7V/5uIpVG6iZFdz
X+qhbV+eAxdYmxP+EpG0uR7H+d6AmNVlVW1tQ1eZTxoj+oNKGARKbteRgr15YMaR
lY+XAxIu/oYWOGC0ohlnc5V3WVyoz9rV0k3pXXzzHgegnldXc+Vgps4mjinpJ75L
TqF/yBE72p9oHTRfQMsOn/IR56zlH/xY6nlITN7hldBfNPc/eCF5Xv7IMn9PP+7B
tF8MFRoF+K1YesjDG7FEtUC7nVyF8S6X9C2z++AoggfrqUqM9xz1RFO2Cx1oqpMo
8blvQGLreBauzyFd9BrETUJ/IcPq6UFVZ9ZvVOpjzTSBLFopkU/n6Q9IIC7biaaV
7/p6LfTd8E6Uu0d9t/EhIzK5UqbM8OvEVUSkXytsUWvH8Pp0bX4sSigNvXbB/3mb
s1SIDa7ToI3lyGXAUkjnLwRroq9UbMYqtuavUSjth4CNOyANlBSQh/RONj8ozovw
1qpoSLAVjCrl61l2eFX3o1Xlr5l0b/PG/S6BGDID5JVriXhBZ7RShVoaHYZIPQLQ
QsUn6tPR9uTUzu418qAP1gMhkQs8/TIYci8fLEUtk1wTQsaSbqnUZhW995nUO3v3
2vr7eYcCHyE4xv57W8bO+ByQ+fR19uLcpVZx1bqGHxXGecPBgrkKFVQ/DNgHVhTH
1nvfGyzJk15rVgAb1og4DGwHmKszltX8amYGH0tkZdQDJTFazD3Mp9rZoGMkKczz
q3GRwnfeZlANQFODY9mX9gV+BTUBpxEEz/kdhOQb6Al6eUb22EEcrUqcSlbNF1Nx
5qqJgTXeIgOPv0X1X+dPkWQsyKkaWP6DGaJpqgFiIFU/GbjZY812aW0JiHru7agd
WPlLJQHWwCFsdJfICks86P/HLWf7f1hbVv3ZJux2TsuRBGKawoQUUljQoz6rKJOR
MMQp7zveTwoqElHm9FTkeqhCjFdfxih5PmfXWGoI0VY5DbzjufIYa7BgkKUYzp5t
YU7LV8C/hJHIrhpxPWNuvT4es9xEsCg4M+R2pYGi6/rxSF9/E7/NAhhBmLIgNwh4
54IYA5opJ2OsweQVLZHzM7FFpfSs9405SVYQ7ImX16WQVmPX3AtnLI/3apeqB1G5
QO3Aw7NX7mt/ieLbYnIwHudEydKoEEBDcJmn0FZNqHR+uSbzByX+MXQmiv0K8Jzz
8VCkn7XQ+QKXC7KVvT7QhgIVGFaNKvneAjm/5hSLYdllTC9sIhm6EguMMWlul+Rc
hxBljbdMI8IEkATX05h/fKPJbL6a508lYyiykq7bOe8om7rv0FDHjFr7I+rkAQyf
c85TVv/7dSKbG0Jlb/n2XD2Zov9s6zH0dhALwueFk6piYceQ0IQyOjbRaR3tOZxS
u7TUqXWTah9a72mYDJ0d4U0rDyvCgTeRkvTbP/aYrtkh0lBnD74fbLTZlPDPc/MJ
ZTCvvWSRYg4mrr9jtPcBWqILB0JlUDHr6+UBgfjUcIlL6jRvSXHvsnmuBB/6xRSu
4LRka8GWSlSVRvzgqB1GKIDq9I6ZeotCh3jntH3d5suMZV1+s3P1LAuXbZaEXre2
WtXwtpBsTdcJrDSUkgjbz6NnezMgFrZOahJquZrMvghE5iSVXRrw47lCA/x7DJY+
57M6j+zIwS+aox3rxhjr7GdV/peM//qMW5v9K1KD3/vltwt7/wMg4xQ9VEYOvcCD
dBZ5CDcE0HxhFkxBaBcpykWX5DQkxvjjSGZYSfl2Qd1iCm80fUahY+RIFOuK/LHQ
QUPEYXX8PlMRKkfQbLsFCXEB7/53IqZCKLes7Oe4Bxo84/9tHbYPTqzyans8LSu6
mKO6DUkKkXtk7zpSRLlo/O1Bv4VtW20qxh3Zwu9Sf47Lf6Xvbnpw7tMHeFmcIbHH
2iHqrXtPicIjWZI3sWlup1AqV1J4GeiltgUkJRNxcwRDl8iuBMIBUT/33Tqx47Lg
B9obolNawIl9HfEY1BKYzdyW3CXS+wEr2qjfUb+xE9hY8NjZvwTERn87V1eoav1X
heD77nj8MBWGuBT8q9tCn83lPKIjK2UNzQlIdOLmRYUAlhjGL6Y5wbcbUWQZQV22
fJC0N5l0a45iaSeOPHE9zw0Yy4IAR4pi4pneD4nHaJz8UqkyKviLgG8EBcROVW15
qgd5Th2d7rGxAKYrOn53Jv4V8tUKAI6QYimowko0Km1gASnMnSfvKHiXILaW084X
6Bro35O0QYCl1vnlAfaUUnc60ldwGEiZRVrEdukSRii3myLXfNviUwyM3Ig9fCWo
xl2mUo85xcLKWL4sDQeonDe88XVFnrThi3OHG+Sp3aSEJI4C3YIMCI6n+b2k+TYt
TkrCnaQ16tbffmWXHlsk2UqD+Vuo8gQd0G8i8RjUCPD3iTKPJexeBjUNBbhKGIpP
8mFc+BukJMnmtJYCzyMOFdNtErKXCCaJMsQ2qRF1LpH33v/+hVP4ZaNjIweg0efj
eb3fHq/DEDKeQtxtgWiDxL/xRNesxOka0X6m2KwEJ07XyxyNIE5gss/1u5vjNqSq
8gI0LRO4//bAclz0wRRMtmmtavNJgJCk68ZOfPI0QeBTZHovynOT5ttQ0mOJOlty
9xqK4DGZ/kizcVpDwlBPtiKxwUDEJwuT0zOjuJP6zHSriOxq4mkXZKbLY/G1n0wf
Mr2dEcCN5pLTHJE6apcDa3XNfS/zRx7xmr4Xf2CswOPSpkaSPdYZt9DPT3RbXhlM
o0TDRnJcNP84A5ASd0DXkVHfB1z/Bf1DpKNgP9sxfq5BEptd+6xyG0MgxWGuSksT
WLEAOmD5IgpwlmUvcbO2tAWCKRbSmfnXHEstAyX9hf5kgM22wBTLR5GA4YIdQilL
5UJ51YEwhNm6sWQJMJdaZk1Kl2fEwcwDXc9eZnvPfSIqXUWgk36dyv9X8hLxVbYJ
NzXUUtEvXUhwrcg3riQDIbiAQHc6tFnSliNFDJKvFPDY/ISZVIFHzvYi580yZnPo
A1nsQZt1vI0Bla2lRqahiJiel2TZ9/xY291PEAmu7BDEVa+FaYwdSaRJascYq3gN
fJJg53vw32sUPCLmpASYH4k8nugOzLuG0g0+8cAXxdXPHMj+dOVYs3tUwFFDa4wv
GHUw4dypDxsrhsds7P9bRw+7kwf/zqO1aD/Zbw6Kfe3EuqgYRG8DAmMn/PsLjbM/
UMojUzn/+QqQeaSkIfFpM4Ljbk3NTQ10kRe3sm0YPLgPDFtX14iPg6feGEo+9L1L
k27XwD1ArIFOvuwu+3VYQdiraHMbDEw/Pfj1sjlfpotWrGMdWsErBStTHy3nIn8w
JJ6MGs7/BGu5mGupW0OEVeGtEj3G7eKpjvT18Fc0AQDFgmcpZW6S9pe+HhXMqeZ2
6ZJoWp16wzIzxcQOSDxxTQlJmpI1NZ5A5GFR2zzyM5lvIlGhrCjk1OU+2JxSQQJ8
tIncd2IX+aTDPHETH0L/0AbNKm1JbVkkbjwc7qktVcDKDuzgTpnzuMBzFxYf2F7u
i41BERBjdY3012zJF1JCXle9JuLMkFN5hp7bjUP1raeajqjrUM4Zr0RL4Rdae1Fx
G+hm27tB9C+0eZpwFW4TtYOrMLaQbDpfjDRbEGcKoR0b0eeRJstjaIsmx1UKzIeW
OWBXuYos/nkyG6aFOZ9P+0NWNbWuuQJumJq8JJGrqmEuu5ZtOxi/TlxLX3EmQn8z
js4tPgRI0rWtVskcQ//oLcgwratqQAsCZ1Zl4dLmJMH7b85PPl5YMP1R3svA9N4P
igVruopG1xg8Br2HeEz4ZZC+5JfCFefDvydaZ+ayVPvUHhocXwA0i+nQd0PgBN2h
kyO0mnIGtK6B+3fHPOVtE/K/yhHlxtbf3NRPmX//p1IXTyxkpaj44w7sOHGvn+lK
P1ZBsijOqxX+aXjAaBOYwEf4+heYsFVM7dbOa+AdXggMWU9hpFv6QIaZfu1CDX6U
fStMJHH3YRZmU2NsxPsgJEn07AZrp3O9aMxIeNAdLOj779Ty+BPRQS8b9D7GXQUA
xxRcdSoRmQjMKOUhZuKmj8QwGuuLuSTLvDWBZsMzZnCVoZzR7dLPGxS+cpYR8nJ5
O1mnYbMufjr3wTAyufOoZ4kdk9ltLNwStFi4/PzkCdisxvIH1XIp4ks7KDmyQ0L5
3FFhjtdTYuQCPTYDTxR6zH7KBi0yUrhsUGzzeKFfQBm6Kv/lYaP08oNKlEeM3wzv
dx7CVabYJLeQpABTkGq1Yg0DV4GKHXmwdB7LUQIwUtPg/lWBWQ4Q5Ve43ZgakqEN
RdUpU/m1rBKrwADe9JfFnEwun+06bPpJr3Shi6n+sClNmXOXRrOCorG2LvAtAwI+
WySN0uLz1kyDysRBCelloJh8p433KzeeRRw4zxcn3uuGEyGMHkiLJv/Yp05STM7b
gYYtuG2nTiR8Kmx0li1TGIc5ZpexikMpb+BIKJ5+hBnVJLhnheKwDo/Y8NotC0Li
U81AKviEk+zpRuZxB9rq+KqGIN4/+/JLxrlf+ZA6jjxpR1dpF3os1kv/VNpzF3xS
qkXLGlULMGizB8jVLiH/vWLod7vC3b5orl6z5/JFxm6+mUJAJgHq/p4Bkru1J00l
Cj9DByn8Epz2wEKZvSlYX+r1E3fSVOUT18PBFpnA5blHGwceZfv4gqhGtvLE/LW9
BL/SvEWvYR6eEA1S/gRY6FeMocGhSWeRWw3BdS/IYjDHewWao3bival2nQQLGJQr
S+Svi0y6E0CCqZGH3CJkwhSQ78gv70rAFNKIK59OuNMNfoVeA/XctnPNcA3YmH6h
0jyum9X+sDzeYhVuNnKpOYPr2f+xPoeew3P9Q7imbuDcm9BvnS2vmlieRZBGuIZv
qSfGFIvCuBrKE1FRAQz7b2SLU6TmQ/JyXycXfgpgZi7X9p6akS0ZxelYlwpMYZtZ
o4L2cpLgu3Y0mDXTghgTc5GIdOmBbjgbGR4XRvh4uExa2rUvikuhg1WU2DIZ3Htt
4cdm/anoXUxMa3VasKXPbvX6ipQWp/Xti90EBubgGxLur1ST5P/zjDM1ioL5xGqq
YcCkWJzKDuNIiy6emvLDnV1AKkgrSmXF1gmYma8BPbRye1tiIz8lt4EbzWgWGBec
eDAHOneG8TN5X0FLCK+kh1Cia7fSsfELTNeQBCYkBexS7bLsvdo89pAdtZLySaYA
Li2pKTUb5V3bKL0yfxp9zFiUDgEVGci4iBS2kGtYqScDkXyDz7B/wMbbCt25Esen
3qyOa2WPapus9+sjorqO9K3TwYFVGQlu5tthrHd/if6R1tCh1UyAZIF+XWHQ5AZE
AZwpke1gXmhb1xY6FtODpYIMGykkdCJudNWSMI2ZLRJDvIBtnGOj0y5mAAGJj1Wh
dbbuBfDb7Zgu2FR5gDuDE0aw3tPG1lF8E4ED5HpoWtfeRJ36GPqru1R44Q6nPA+y
BF6D6EbWEEIRkT7eeuDY0fDNT0pJdTQcIsbOxcqtcU765y/E2lXXNP0/2XnkKLGJ
h4ongR3uqHSaAHm9JoFpi1VxeeM1QD23h/YCLWmBqSBaHpXtFAQl+dNf+9zzytl/
XGPDI/tfbDKgvzBiQppft/w+9qzI0hj/c8xwmwj8Z2firJyaTSGV1JIkzJquWaAN
qGZAtQ+H0d4iJNf4ZLuCZOO8U7xsfyqMp6pl/+r6JuOrtcF/gghWKStXSw5Rm1Y3
EVv9viWNpH6khoHRrqoDWMflPnnzHJ7xbC11ztpHgnhBJXVdotpcAhMutu9WUxSd
C5cjtQfhttvlUQrNdaer8K5B1FyD3WJtK9yVeqEQAGYGBvwv8qudSWd22fqukK7T
M/n92DDM/xvwsNJVml096LjkSaTmv8cuhNfrSLCX3x1Z9E0TElovdTr3waFPqYMJ
fPo1wl3VpzYeAs7K3BvN3u9JDLsEdnz5N6X1ZwhA3kFuN3tUhUiKNn6WnkAV65Ks
WM7ex9+kEMeljd4f7stEDqeHZW7H4pjqr4DfzbVQt/7+RdfWyTZatMEoFoODAavs
L3cwSVwTN06b5wesSt4i9oy2xI+d0gudbonINKo9yxgWF9vM3jzm8GsDwG/mj+F0
T0BIxVbCIjsvd+p/0kXWIVZf+rl8RWRUqrwQFFWJabRIy7ydxZ9CLpGGtskj8/nv
voG9zlAv9XqX90Bu57makr+/+Lra5Ood67rnhBHE0nrrmmJN1LZ2haVc6xhbarEb
j5sVFlvnzlz9WdeIn6R70TnerSC2y+AfUc3xP/Z9SyprmaKlfDVTLAyEe8hCqZDZ
k+s/kxTBsXK5XlfSRL/WOBkkfs/ZUlL9zAA1NB5+NvOMd/xvAHeSonbKd+Gs5AI8
OXrofNLid1TkibvdmVKJADyicH3KeT/S02MIfWcX/NVzwxR+fMPeVZpUmMsXkOV5
r05csWrAB4NNiaVFTVnXKCnLdsc2GPjazbzROmDN+p3uRoo0O/q185+joFDTDgWr
iBzfcLXDnpzT141c2fMfRppLDEHEvne+VHRXdYSOjfUdLyTW6EDs/nynKH59heqF
RhLUNAaZPRCyKO6+tb0oTmg4tlzyFIC0KdL2FJF8PWNTe8NWmVyGusGux/3SFzzZ
/OasSVJ7/NK2irRzzdsauzzIDSOmX5oy5UOroCxERKoSAJuy1899bVeKqdpJmfM0
Z7y3OfWX/LcgP80RU86SBZO+ReIhBxRaZRbe/PELiCvH7XKREfGuC8bZtrTe/ATE
ffaCpn8hCkfp4JYL5DxVv3TaWiJq0+ftTryx3ohdtG2eKOCukdQdUm34q4Y6GaW7
cXsjb2DPvS3LqJvpssuStSXVpnNCnWvTis2P8QOSoeC+3ZlxLCyFuwkD3B1g7ga7
AabMo1gOlHTQZJFpesLtLILjt4eddXXv8cdv+DvDpmYq2tL7Wb20ARvXBHUIXAEc
7QC+Em6a085NsXBoouqLlVvpH6nhUWikhTuh5oq8FKrpSdgIJ8tXGF8Tzy8geip+
eO2xfdsfnYxBdUE6NMXImxYfZTA8l4TM34faFqJiPVVydNX1/79/PrXPuzZ2WdPu
U0ncHvS31ho/G/YBwrKx5GHKdzXFlo/Io02U45NScrqnfW3WgV4fHOt1WBh2JH8Q
MoLYDYWta6h6cQKwfmhdGTKar7F67w5J2ub9slHaRp269yhuq/9btJ1+U6NxSI10
wExiMTWiKn/NWktunH7gIO9KCnA7P56a0ZrlTsZ+c8XqVArxWwlYGGkMPJbZfcDG
9vWI8VTjeZEHJ4xLQOyp//2Ssle2/NBtTt9gub7xvqa2rVLIcyOA+h4YwcSswLyQ
Nai/mTHRtp9SrDjM77dYHzKEU9LBHA6mDqPDATPgSDxkc8NZISoTSJmzzMCmEukr
2PjuQn6kbEMZFLz2g1JGEbMCg+/Uh2kII2bdWKQELIoD3BCrvOb8k+YSvqB00MyL
d2syGUFjRvFj7MchF5QlOQrFgroII/iqWJGSF6S9/bMwYOSC6yIG6fmI9vsVb3p8
j/8HkeSBnz/NeGDz8loeS6tiZcYXMsFlROQbmBVMX3Mn2MZ7Z5PIA7w9caNLTllJ
WIZt3ar75793NiHqtoLAffPztX5o59L0RyGSNp/zmesMpn/iZlqtWzRPX7D7tdjf
BOmvNrqHQk2guDrJHblJJoVkNWeQs6Oshg4HX8Ir9t5+h+QnYA7L/Hd3uA127/sQ
gZOQBM80FK9Nib+rDipBwjNq+OHG/Kq2aleUPkmkLnby4Ky+rNizz1Sf1WiMhmzv
fWsNqN8kzq4kH+3cl3fqy6efaW0MtpPpjixu9eCxiZS66Zzh7X6uQ0b0QmJinTxV
GPaCGsRzd/0pfpLnH9kohIkVXWaCQfww7XkuRa2b6alg+mBPola6hCj3EwvKC0D4
mQJ9y6hY7Yl2lJNOenajjxbRkR8TdpBQGy0mUxsdGb+Zbp0P9ftSqfIus7D449s3
O6jKoxQB/lkBpaYSYxhoPuOguHo/X7z6TT6y6KPA/gV2gr9sIRb6Ahd4VjwqXO9l
tnfCxq7M13UM/WDkSH/lQmkZFEyzw2xM4b2yBjjcF/9h6fe2XepUIFquPOmhiRji
IXu34RUyAX3clL1xaQTJj73LLi498eaWFQFacnbkH7LMxfvAp5VVW+1QDbw9vvo1
7C7GCtAF4nXclpy93SdBJXLVzj/I6anxR6lQA7ViZ3neTPfMkznGHQndyRqtXApy
rtS1CsKrdFIMAhWWRrCpjguKp5CbBngRh3i6MzmxG/g8W0Q+kLMR78hp51Y5mfCG
+qiO1yTrF//Fmk7IdFU4VDFW+hqeG0yOwFGVucFExeNzI7XrP8Hf2R8cbcBf3yWc
M+NUyvFSJwQ2yAkFn5ctGiczNt9KaRHXtdjXob3msZVoDMYFHRDKXplgkXRZMS31
gQVR8VE70ud74ZGP4WqAHJhhg7tyzj4XpnHspVwo53RGM1rdWtuW73koAqV5X6/d
tE5AYj+Y4W4OVpPiGGq4sOUP+heRfHgufd/oDR7t0zyBlk+WO1AKC5whs1dniMNE
xsJsSwRqg3nIUkgZHNvhFSQD+v3jxTWusjQw9suwGHAtuzqKwF2PnC1CAL+0+ZXj
ET44sUCf/U6pbvKakHCo4fFrVtVcnXOFdKw3TcdD5cYXTDOhYzNXXBdV5cWBOMCv
ZA7lxdh4mWwPNmwBT67xwUVHI2+zwe5OJj12odSBwcqEC4oEX/HtmZCX9TVbaqw/
nDlOHRk80neDEaRLIabxZ0azaCejRoWWTq8jK36p3nFBjecQMM5DTfUecJ38a1F8
Tt+P+jWcdnLI9bi/f+PSMTOh0+tmj1scel30GJ7evyUmnnWEB0WX8DpPP31gpy4U
+eg53kKh0YolSfGn9AX9vGq12IfFjcNx4cJjRhFOXhh0fGoYkPEviQvDb8hAF5me
t777FmPwB6F8ZLET7xPEqN+F8b7dql5TJ7LQH39okXGbsGZiF1fdKC3tJizhrTbE
RHQQ/QIE1G/M0FkKv4VUvP0moyQUEAF/KaSSjVeAEwtCad3fGxjN2GIFeLc80Xls
oMk19/EF2FF+ZwwMcnVdLwiknxbEbqvlrp/d4n4IDYaLlgYo8OR0ziyU2KAaLODN
CXt9mf2luWf4o9XGbYo66AIcZ7Y9hyR3VaIP1jtmt2Ba2Lq7gB1pzLSquIJV+eh7
qQR313PTk05Xgg96kCEBtY+gLDZ7qvi3qX5yDnMptKdBDH82jZuUuAbbcF7dU047
VlCHDvJN8XC4aMobAQfQEisE1UTgfEwp0VfbB4sA3abIXezbeTHNGbdbXt34Rxnu
3fn+Hm8XbBRUJA2VCz6IHv0ts9Z9JphoNbY9LpORZFvgedvETo2g5ADBMvS7XMRY
y5sOGcT3Z3FfLrwxT8iiAdrlr1odQ2pOxM/hkUPyLCoz5t5AkExNSizwS1ix4Uxc
U5RZPBsZi+vqzqwFRL3nHJk15YwRl44U+pG7UQPSpK3DAWiWfRIPvbVNhnu4MOgm
WsZL+iXN8I4Qm7bfhtirUsE2qYa9vdzhDzqXTfvcyTAtVBE5fgfDnoZxdfhNrcBr
2M0bdC6kOyTVGO+mhCO7R2wtPpqDioTha77lqklRA8cLBnQ89ZFj9BgOxXF46J72
1HpCz5zdArkhMoLPKQKWjXKJu4Jw7RGnx7WPQILMguMPLXyn8QclBj4GAGh+LogD
Vm/J7Uy9fDbpw7hY41XCT5jFG0jcTsMBatu5XeL8rY+EzFh6riQ/gKIEPOm/dVJE
Z2Lkvf0fB83EuCrGw4xeEXCJcRp+T7c2sV4Evy14SVf+OjfA7W99JXxHgPI4Qvf+
kLmJJXrOR2wBUkPcUqZVNrMndvDxRdL6T11r84Z+T8bnDre4DT8VnqSH+2YDXe5O
d+JvkYlqUv0q1s5hOGGU0NOPqFoY0mdfueieltYj3RD8qODcZqo+1YKDqKG8eXft
rG1IF/O+2CmBYxksPQLKSLa6WFtQ83PL2jKb8Q6J300joTSySQGrPNLRedc9weDe
nLj3Ov+Ooy8p8ngx5cxb9JNyx/PUebH3wQWNKgoCBUtXneJ/rjOfJeWDXZHYktCk
ep6zYjGxiLRea+6ZvLT7ac9oWkst3X6TMuSsg2rGLxZPuvORW3FLE7Qh5HLlttIl
BjhIFsXMY4zpeImcL6lTDKOztOV0JBo+fjyoINF7XJf4G2KzlPkA/OlR84kpGD6v
AGYG0XenBuLYSTsWSNcPMkXPf3G5Ai3EODxWCyyuhamqblxFV3sZUKhO8s+eCty8
EnuWw0SoCw4bh/CR+LCCCncyyfz2j0y/U7nFfegt6uKth7iyIx9d0jACAA0epYPe
7jZG+hPcJIJwX2/5ZQGAF4+9t8JEWOqdgA/HDSuui+Pp1DxFO006jnJSKRkav+Fu
0jGPNCbe8e2XOv/ydmuqqA8IFJqp9ukaXZdheMIGtdJ3A3cXh9RmvKlCL4sWVLKS
+Jl/lXRlKkGm5Bh4Zm5PE3oyHGm74zNOc0VLcNYPxLItReQd3UokQ6hyEQeoG25a
k6ovBLyXcbG7p/TS9zKZAcjmfaMkGiF7dD3VhyqOd4GdXlOsUVlfx+4aH95fWmrJ
bdHKVPxCVcrwbUkTt+JnKJTG5cg2TWL9PAYaWiTMvSij4VS3dX770kVJ9SGJDeR4
DEarQobfd3Ap684JH67EMKnz8zHxRvoGgNgcHaU5ZH3ZBtBg1E7ighJGCVDXMFUz
2qxDxHgQEbCFeVt1cZRhQ2cST4Hzh56nFgasqJ8hGvnytXz0Ia07r3DnnHjv3ulF
/zus8ln7mi+UjFUS/ujIXLdGGNK8egjXDZmheVwvxgOEVCNbIqPnJ3cb34BvLbhz
0mhR7G3ID+PMpI1yPXXQzz7k6sQcEzmNvjE9vwuOFsz0Rj0lgXztVZ1uoRMvQ7G/
6O9cgFlNFrj1+uDCfCwvJ2+TcTx15THZdWDYV6ezasDgfJhxpZW+2o766pXYyRTu
pw3WmiamWljLywmKk1BA9PsXlieOKbyBb36xDQXSkhXRVC+US8C1yddJR04EOzCJ
YI2MBH4u07f3KnsuvO3KokoCooS1FpcGPVlOIhGo6kMhjmNr7E/m9VoLZiDpuKXU
KBCG2zSF27PxgnrPlPDWOdmOUb10XljDPHTw0ScW3ARlGuysIZ4wQhc1JW5GcD/5
YRiA0vdvp+4lO2xelvP1WzfZPQ64pPnVF9HJuYa9BkT7TqZZRntJ1swmwdxFe5dZ
mjnYMWhkzVpW1gSphUvqKOjlCfi5JUHvN/OAFgP9Suvf6fXNEobrVmkatRwZ/5F2
jERPfeSkjNecJorhLgdmkiAyLuLR7FneLfAT76xr+EWSSWg1Y6rIukRNluoPQjFF
gitjZZSkACQ7kkie/Cc5q5Ld87Z8sPllTOT1rzgfnY4KJtzsBtGzATqXp5coCeVE
m2jCL5vgxMjfXsfSoJJobqiwqGRbSA51sC5kkJ5vui0etulCelrAO4/Jaw7yI3rw
7PAGqogfhWedqChG4rqLool2wQ4ERWpkbbpjOYq6CAAoDmeUB5vW85UpCYkh6sXh
s8cO4e8NVFF6JH3kwhUsSF4b8TzbtjUx8LjGtrK2ErJwhoe8l7pZ0C+fz/R1Nb0b
BiMZoKb+XBn7rSNtl4kM+rNIXNujqvJHy9IgmNYQn06iNQHpI0v8oeEGnrbbATUZ
Xr2MtuM6tw+R4YEgr1c7HDrScpU5M65+pThSXd5DxOhvat/wa8t3IedXMt19T3qI
8f/o8o6yH6IlSZrgkTVpmqy02zIWmy+/WH6w9XuEN9rIAW++jJ86Do2AqRVC3it2
pqlAsrQ8+tgwIf/l71+tXadlRRzr4RtBxgXzrfeDlJLcJE5DBRSa+0hK1fpUV7Ke
+a6zny+ACur1Vb7c2EPZIfRYKmPDsNSDoxxyBpors7TZbukNqduLQrYEZKWQh3Jc
ItJvnJHxuWL3bqIuirCKVc34BhzyVboe1fSRYgTlHP6E4l7f//swNL9Q6QDUJhJG
MEdge88BG9cawYRWFWtEbAKNSwadl10YDQdCelKOrkzrZK//tgV4VrKfugU5JaEe
eBF0Icz38cmf5ABiXuoQxEsjkMg2t4ezKEaHTcgXLMrXnjM8xULZ6chHpRZzSWnj
p9r7umKaXs1BCIO5YNXsW7Vlh0wKyXAdNfLOif85gUtiXuKdUHOSjbPhLbmpaZ+G
a6wgbdP/4AylY3oYLofBzY9hu6H8QFjAvFJVchEmxuJsUAyGb5sGuU6Toz/D6hph
Z+KyL7NYyPRRPG3QmWfiTEL7i2c00QsKfwe+xl6GkS93hdMDTbor5ael/84nYLtA
Aj+bWwnOpHX9OU8KLiM3hZa3hOIyVu9cibfyuXrgUk1d4y9UEFSGTRTwkjHGWAea
b+3zrWJYWrHdoO7Q0aYL8sYxQn1rsHoj92PUWHdgjxLwCcwTo5P3WjdfrdE6I1di
iU2+jOULjZLC9BheNklBX8wOkRe2ARoazIIDXRfK/bvLbmoW0+rLDZHK7wgKHSPQ
ipEU/1cJkl5+YGd29YKAWzIbcnV6UftiIGmQAt5WWd9nFNs9NGF/54mGwMUc09fp
44Eun6vGONxCzDo2Yilc9mcXfIccGx+nIevCN701+Dm2TVuotnlAMsvMBmcc3DBG
o5JsvIAWVN5wp6AfQZ/PndOPH2eZtXEhz+haWb97UjAiLy/P0BXr8QjkWFGY10nQ
EVB8VhAIO5ZQAQpzyjjzU+RzPaoPu2FjJwDoJwJmqmSTO24CPm1MocWp5uyPPF+P
/jReOEu5vjCKidvQa3TvvQbpebLUia7oEOzew17enR3xc1kT0ZfFDQHlKDsY8rRV
bkZPlfs2q8ic72r6WlhfiXoGKRyNK1mgXpUEo5dScsJY+6CS8E0jNIRnt2PFS7xl
YeqmEJJWm1FAX8lBSI9+HUOPkosBMtlvrjsPPKGYAy+t4XXpVco84n1hDAxAE9i2
CMiSn8wcBx+Dg9mm5jTwhXKSQfWTb8bcWwtpsfyX4qhDHr/UeEmeqAAZoBAF5lno
jS8O+kdDdUvTYgc3tytv4nu2bmNgnuPgU7HqbBhilCh2CRn7k37gtAlV7JKtapJ+
FyYmWbJeQayitg9UTp5pbvyeo1OTvQd4o5G22Dga893v7EnKfMF9foWsJIVznIJq
CiqGW/Dhw4KK6PtBZld9VXBlGb5C9q3+z4GviOqXp8Nb+DS7oqyjXKhKNCXQeg0f
KOUISu4BfyYFxgLGVlafFKQr0jtVzWtF6uhCQPqobT3h+nQCdXyORQTHAv/9YJWP
2IoA11/9gBlTGUldqoD0K8ndS0QW+VIVbDN2Xeq80EA8nBANg5aL1dTl3p1etU5a
BsS94twoH4cUM9sfReTtNWHcXY57nHRBgxNpES6O44YmhNIzPvHaw/nO7w49B+pB
p7nygU87UsDv2lGznQUYF6jKOtKXMP4b9flyeQSSQZxZMDQDP1jVmJz+GW8bJf9x
u7/UIch8TAFmks/1a7orUrRMYjPFI+ejjJyfZnK+VcRWes2feiT/5HAKCxU06riV
gANzcwyI61w+qBNDAceqmeLwDrQGF21qOh2pDTp1tY2wlJ7uSiWk00mckXjIvUMZ
zaIqC24OpJnnt+AOhSiuwrSves5nBngwisESFNDXvj2ivO0oDqyhKAU8JEOaDpDj
7Z6WBfKV43C1Y12ifbILHlxp1cAWBIMQjENdPIzQRIAkbEobR9ojeJDL5nlDOaXf
hCvNpuJCE9vU4brzUla4ZFw7N7oLNEqBZqEs2p0QsvaNOIalc3xjNATgmTGdH760
y0xC7Mjrji4bZwsREnCAGn1v5hHbMCAlEFqsv8aXP1A28h/hSPT6BP5nTsIQKrla
CWUAw7dIiTG5w7U25XoG5ksVEEi4+X3YundHGs5CONbJmRPmHL6iUKUj7idMdA0V
uwnrMUZ16tOVtTBs5IdW+wsj1XPDgNJAmj+MAl1o1JwXWzm2bNYZZWl2vgVZPA2k
Ev1FCh03nfIQ8z5P8UxQzoYxu1ZES46PrQ4rBj4p5raso0ViNPDZlcv1xd7Uj1s6
hubbjkyV+toGmHng0hl8cwVNXAYscRJODSL6VXOM/kujQO1CGlGJ2cE2hMW2lEEg
gUbp1u/xq708r6qWZWOVYWORZ57NMcw+9DBuYHHcE78YVhQB/Cmbb5uFpdRd69Ew
+i78nOd6TdlJNFhDrCPGOU3gY38FTvG22PjneDQU068GXSthAvyWdECFhAnyNVI/
jASN/ihcBjq4/VhQRqctu0BbvdNoUYqnZeIqn8AQiCMwEwgKAD4v7K8yWR1vNW9F
h8V8oS7PAKkgpVYPF28umxHNKPT5rq57cM0zdygRneQ83a+FP2bT34a7apsjTShQ
3CVH656BopfLZUEPG2/Vme7pZ0uKJV6ZfQHulvo44szgjY017dXP+OVXODpG3hCK
mUb95DeGN+pugIH7yFKBcp+ZRtahHyp+YPMKQaRGMhbLrxQYaNChFx5KUBuppwH6
MZsbDljDVv2moG/4G9j+0epsmdM4K3iEdKZnaT7o9o5gZ4z8nCTl16hfZKaYYT8H
vX9YXV29WJQ2wI38r+wLVHkqlj9ma7vD0EuEpViVHmnlwQhx19njiGSK7gULVbb6
XQdAQ63vuFeU9aVFht0V0NZjvgfBD1lxlgglEOR/DlUEQspsemWSY43h6ZJner4S
EDQqOHFezYItWX7oevBJyyT8b1YMrcR4Hl31h0UI1xxPda16vLZaZxVV2z0/6mlN
RXCxsW7PqXmwxRaKCjDtDZ6WR5VHEEdqCgYNZMZITUOTOhduy0UkgUzoH6sX7w/K
hlmmYjBIyO34gZKL9S2jdbPOZEJUmsz/jzrZ0ocAlmJqVldQqSnz+W7Dyyux8OPL
Rwiov6snJmiLNg+vlFIL1bchqveX1gJ0CL9w8pxxamDO97uH+uEE6nomA/MjR1bj
r1rRqfVDVf9Mo3iwQEHY7ZaWOZ1gMx/NTum8m+cEtemir7MYMOEUpgVSl5zpfpT4
eBbtXIVenlCV7+uEwUV+J+4lpl+98uUr1GPWzKnR8vr0HdTQPX2YdoFzorQfqBGz
HQBfrVR+oWtx4RRci2FQ1MaK4MHQ0YAWTpvzp/lWXamHRVPphaxuJXOKgZcjQl+Y
741uLImKyLjPJbCg1HBcCNiYM3IReHxEdfcxh1aMMwnuyZR4TN3oLw7JBvNBy62g
twBSTTGdu2vqDJMv/4pCvMAo0raQ1bWmWe1qsU5vRyFP+QtGe6Pc1G3af+nkuYuG
do/zXnCHLik/BHXKrQDOrNxWyTGAY9rJVlm8uJPa/oujQTvgAeItIYnBHiw/BfCQ
1tswVZsv7uH/sgmNe+6vDOU3d9RRrmCOrzl+gshUNqOvZiUt2r9k89Vv5LDVLnSk
S0856euoeD2kRnDL4lLRUU3Ub+nxveJYZQe6b4re0PiB7iyv7peKtll/9k0Srtde
I7JggU8Sjk/9lSfLBySULqMMct0mmdByVfwHOQ8VmRFHv3NL3+2wpJki4XcoJWlh
11GpFvSnwwqAr5Zw+OLr2JEXrbhJ7oxoDrDARxH7fSLbrtAIxWIRwXguhdQxWUcy
lrMgXlQC3Ij0VR/5q4sCeALFBS9N9z9kE05ZCLgb5xC5PfgKdWMXXhy/gwk6KNbh
luQ1zfnONXqBPcOK3qvu4lzPLgLp4226/rX/iwu1G5QsgcdyXjnt878ZxjI3gJts
TvYcn7i4XlDmUp3Da3k/5/OxffGNHvmXNAhCEL3JiSAEWTPqTWxDyWPqNioP+Ito
EttCIrJ0alf9DdkuSPVVqco6beT2mLBjny8Gw5kU6VAX9o57OvXlPjyW/JylI4Ft
m4LqjDMUihaYMz+nSt3FkgKYaBzU0N2mn3ikvnTvSSsb5Q9UIZpP6yuC3e3nLqwL
1k/V0mevhYrmnfdtHJIbwBFoqoFupeRh6GCueOKWYlyCuwhO1fYVOGmZAQ93S2vj
1Xgd1wCEXwzfaoD51ehSFSD89nGegc4lbl+h+Nz9biCqMNzffqe8Q8FNfspBN2Sj
FGZ1wV/LHd1jC/kg19jRdTkizLEWiRKfc2qaqDHxGRRmCUemnfQqaoUKGgrI3TCg
vGW8uo3gqCY4vITlwx7wl+/tTkQRq9VBdNtcr/bTk/QkaBuFQZAupw5QiMi+cn7i
zFz31hZk+EvyI9IhlQ5pt4RL8xTer8BN2h9viHWFdLPDlkA3lZMUzTIl1MD7rY9i
XIm+sQxATp+xhJ8AAh7rJNowl0KchzfECerkpxoRrxhXxd+ALffClZVvo8DETjyg
34cCp1VFqurKIPFKnQ5yNFMEnYDMU4vrYstt1zIh240fzBjXfk04cm9L2WfysAOq
1K0o0SuU95Tdmb3DoLcs4EGNSelzK8KgPD7C3u3v8kLJXCoK43zit2VUKWKoawbT
j8s5QN6FgQYr5228eO24iZF3V0KCgQ/fvMTgVTXUrzdMtX/EYy9am9LsVdI69WiU
EdpJ7Fz8CGlQt58WNIWODqwxImbmo0YdrUGuzAPuFii/mxLSit3bgr//WreJ1wRo
iQ/5Ms4scNW75YRy2lUVQ31O7HG5wYfxGCLbTune3BGRIL5k/t/oGaGfB5YXCdok
fQRewQ1DGUboW4NfnMpGurNBui07SankuTwP1KvWu3d6HFM80hY2gdf5lmyeQgmM
beFoUSGwX8enozxTl2ciijLc1IUaSd/TzkIpW3cOUXnvfd9W1GNSdYuguUT4Dqnw
fJbHhMtLkvASZ1+7L/oLQDpK4/kqHdoLjFtES3Hj0H5BZwoJzrxZd3Nih9zOJj1v
lU5S+QRFsBEZ1rEZ0mnPTmolQnnXn8lIOQuGT6iGxSNExtPzOaYCnMnkmjRM/KvM
cKudXSNUrXy30szYuFqVTA7ZNWMuhMSqGv95p7v/cp9qQNzljlj5rgmmlsFI9t8d
QeBqkj+R8r3LReDwnB2OlAyeo9z9HlKK29nvV/l4mNr6A3QCu5HDTvIWVP1T8wOA
ks2AMASd0zfeLLMEu1iqnsjM8JsTjt1SZRiF0V9w6i7j0WYyIAtY+s/3ZRv0rgdh
oarf8pUK3Re3nbWwfScZIO+2pUI3Bw3E2eIoFR8WxCvCWy3aLvRAV7lHfcd9YMXC
fCS9gWAv3uwBBRqw3EWlS7w+yDB1NinhRSPWv/pdhggtrKV9MWSYIubSIWY4R+tH
zVn9gknauq3DLqA1GxkDmXxkQzKbSgFhZqiiX0wmWcAzWxQOnw++F2pN91m8y5wX
USMAZHobuynTHOYXR0E+X48Ed4Hc4Z0zzKZYTpE2cfvUm3NASgqRPkj9N9Mw5qgt
MStcJRvaZ58z4JkVkds4bzRkzQVQmt3knIBhEhqRxnYLioDhVGZWvQ+8Q1Q+nU0w
FtH/jqfHwuD08E/wZCOowR8FusRnB9k9ZPHO30bYlc8XSlsE/9ASmmy00iXnq2PD
LQdmN8wW+PeIuz9dajSp6ScrjXmX8dEg590y4iZMhDUcsVn8zVKMkRhDHd2ZTRXL
4WSh8rQ9RlwVZolWb6JGZEilQqIpKXNzluZqWJxMEL7HVLAEIap0rylhyBWuWmQ+
mr8qkqcKg2xpld8PvkqULVinrSOc37XuUkMs1DMqTdbio0rqF/QZDUsLj2KOhEdd
z5CXeEydiW6D2vHQyn5nPDIo0Z6yGOzAanbYrRCcZyGxEoK/wooKz7HCv+jZmD2j
Ot3uRCunvw1CU3kdifSHZZhngNbJSPktqjFzrvK8eKbOI2rtQPPh2SpmQscuwWUk
lDgoVkePcqeesW4pBBj9+sVgjwF8CPU27O0pZnifVf58cBTLg2Ho1fSfAvUTOSAF
/Woke+ubHS8+KeQ7U8B9TShJOoxqTO+v2m3vhztKpK+ZG9KTP9BMW6f4BA1me0w3
AJVwG0mq9KtZTyTrRdDZPWVJBzDPGCKR+zAwGHJsNfVkqFORwnogubN49dXurk8X
JCiICaoZPJKK071juTCaZcF+hXYnstKym91U8+AEjy9kC5b+gohvuKIF5Bc9RCrA
iiViyROwhPrxd3YQ4XfatkKN/jN9GwKEWnd9rf+tAt3wyBjN/0sUtU97yAezbkPc
HY7rVFEzY4CJ+CLztdPseX3jTIXu8MZWh7TiOY5/7NhKu437aQD4DMKEFfzOEC+q
MsGeg68YkMFH3xh5RLuRRT7wWJ4qZDH/+B7w79ofgjV9G1eGdf4Ez8YpslnBYSS9
zMQN7U/YAeryKT1hNXtEKRQWDT3LlbzVEdxrZhiLBDekmxNCR9/J7Jm0GfCap7zP
NdCy3BS5FwslmXYbWi83/idd3Vu2A4be1EH6XS34siXgHgsM27s5cqQTGTuvTrWJ
x77RaJB0WIf8AJ/WzEX+JvgZNkIAMUCuJRPFc1+hUMAZ4PhXtdvvauHJYnT7V8bX
67bFDWVsSCBgxtLKHMfTz2yUan63htHQq605RHDSW8OVWIXFxEUhjk9fp8Agc6MH
TkFum8I0EDadGygxg54alNQPa1ZVR9sDflin/jMKe21ZKS4S0U79mmfhUm6zkhBs
aWNzdSNfDBye1b8dJqBMLAPmz0t4p3fidh5hKxrBnqvd5H9BQrPcjGs3KOAoHHXZ
qF4eHVERACKfSjO8EnWvYhfR/iHOqw4jPR87zoRWBMD4es9ZYCJchmgDteDJT8DK
I2hJSZEQh5Zc3AptCvMZZ/8F5VebytdP1733FAK5PjrIFXQh4LJ0VDM+nPg8rz40
Bubo6hUiB4DrmOSdSetlcc90Ylp6OySOBD2Xnz+iJv0fT1k3Qd/XI+9d2xldSmcI
Sk0MatQKtPCB0FwNNYKyTx4FiP7bc6nRhw07sp9+Yx27XwQP4166FWM9cIM9CHpk
cs8QIZBoMx9zi5GnhCGQxRNQ45v8Fvfe9ctuk9+WQ1PYmPxavcNqCZs7FNzqC8yt
L6V3WdyK35Kqasj9vaaAxt0Ch8IL+IuPFoeXWYd6Kw+qa9OM0FNUVyzUjNS3DDFH
xMKttGRITTx33TRJ0qjo99AEfoUWZmrG+aU9pYTcziekurf7yCo5Oe9snBBu1A0H
tmB06h8NoWrUvW6WEbdmQRECyIgpbHURojEIU8MMEyioUz+JD+oFgveul0IAY2ot
NBD23ZI6nOrPMJndq7IbgVhpSHRb2+zlqUdpIFdTN20CupLzHD79Fiu0rCb2g1Dt
TKzjHf11YuTKxpl7JDLmPUWEJfnB7yahgq+ET4GE4N9itLdkrtrU60NE70WgbZHq
VuBJupLyuXeZRWH4Oto7HmFfiQbRfeXahfDkRzRcewsPyRNHWP75oSe/B/WChpzJ
ejufSeAsnyeVZgDs3rIju7LuuYqzJ19n+iWvSYPXdo/Gi3PEjZqtXq2PumKNkeVY
Cyj0Gx6omiFNz0zwpZllXJQY6yoiSqvWqiQEJAmUv0WP0vCNjfMk7a1fXh03S0bI
tel6JMS4bFM8kMw/gz966GIzmaYi2nkk8i4fys9cO1ZRT2a5tB9mRVySv6w75OQi
m4c/4+eJwXXQOT1NRa+9esyc5Qg9RMzkdcE0ApdjDZsAn3O0mAbOb1UZ5LO32uDs
hBlTjr+vA5GXRDkm+bxoaVfbTO5hrHnpwVZj9dOxGr/Xf0IQ2HohSkb5v3nnkyeW
kNEKOW4V6UBsuzV5C7ela9khzn9vKv/6VKiI2fzKwjdHxBeR9NucD88m5SlzLc0w
4Jr1F1macmQi/f5jSUS7FpFYYZD7zDjGOiV+RnOJmNtCeSdjv9dqt7VfLPk7nINZ
fFBDqDJl+WG9+QoLl4QcWArCkkeXbIF0TLlJ+C3/3erh8MXzp5zUs8QV2eby5Q2f
D49NBKWDJraB4FRxOj9Cz4kgW/m/EG70506Vof4xrB4knlpkwJGrxtPY3dGNznai
+nNq0YSDu+nXc2LoHahtLsa8Hrf3Ehx1qRTwG5uJZyXYmQ6hCy7m3WG1Je8bIWS8
tCq20lJse4En9j5IoP36QCg7toJPZ/UN/kFQH6WgBz4tUMXj5gxOGG+j/3Y07qAS
jaXCxNG5XKU3s9SalcnP4B3BgIeb9zpTAqCKaRMHcY+x7brdbHF92PBujQyiSER2
rmXqIFnQyLo+ZEUkeOgwh+djSEYLuoQmH9HswyBCCLbsrWgqc6Brhm4KvoKE8Elj
PeI2/VNly9v+tZjUty8Yi1MkgtK6BKUObuV+tpxTNSFuPmFVCRJNTlprY7LeoGX1
udVOxb9MjEl8VfSa/78iA50kFxH5B+OmBHvIEHkxT4Ch0W+e4H99ozfd+zCmfL4n
puPw3RYKI0fEZIwPP8zKyrq3poBI6cg+1p+p1u33cCndY03+r++8EFLAvaAkiBmE
P3/wCPC+7SJHUyLEC2TZGFMoCDKEI0znvyx+xFDTdPNIs3BgPr0WTdg6j03PxJuO
KfNIacdr396mec0ySQ2YvxOtPqSvHm+HgXMF81MwTbJs5/HwKs9J4kBXEHdxiyyw
VzMUz0fJ6oGbz5CIbBw9ZnPW4GyRMRqrDWuvF52mezXhRL2LoLcWrIOXNFhnwYo6
GVg4sb5J8rGVptcmABCquzEbjS1Yy3y58VxAJsQaBmPleg1u90tPusHOZsW3/04X
okGVOvTGdXNUqWTVmfxkxeb5eqMAYx/Q7yaGz6xHHX3DYa8/qHGCbTYQ/UnU/cbz
ZWT9+dcxbfX7QgntZhBMaCJot1pya1CHWZ6ami6EV/vSmmWjCSkFaQOG1fsa8Ue0
3cFjizRjLW50SVBs2XrAfXLgDb5V+UH04Iu6fa60sJmHqZ2Ffu0nTAMQIdFwrsXP
s4t4+Y0VzrJ3pxv8NN6F/aNJI9WOz7ivdVu5aV2yo4IZILZ3uHtCE2ajg9V7Ph1r
/yXRBk8OeLT5r9Z9XC+VniKX+RQ9FYdwzw4Qom2p2ISB0PpOoEctN+n7WmQ4XTlf
WFN5hoArgK+dswsuaAdLCqjoTtwaaWwZpMTU21E8c86aem/DjsvUeKlG9JZcvEO6
JS6BiX6sXNeokSiGglx+ysojP50Mc6Q0IRotDln/ynBTfs0XGAf/hK6+3IRm6N56
+dG7SiL1q4AFiibUdpgNtI9ytxYTbCKMeVZQ3vtt6CyPGWAhlJAxljluLyzXuK9u
jDWbXr93W+/S0cNXvmbt6HS5XkANJPxSyf855eXTPF7BaM1F7WPxAuQ/u/T5jaRq
6DaPVfZrMQKmb/7T7EbE78BNXI9lvHeVynUPxzd6lcYv7k4dbk02eB0QElUoGX3Q
aNpFYZIxZS2wsdIeE48+0th9WaIVGtzRx1l+oQDlcR30G64gbO63ctUc1vegGGYy
/CcL9GHkUrE4hhTGcQGIFBE3dP5dkwg9Vax1b0t1De8vdmJNZhG6GcUlmejumQai
hjuCqRQWs60yvb1zbeSNNdxaI8j52Vc6uuixSsHUIhRBRqgS7d4Zjb4/KvMDXUVF
oMoU2frpnZXxlp82WvXRKZWZvP41H8cb2P7MxsDKOpHvoVYd4r7IrCExYYxH4Js0
8nn7kmdutcBKF3ruzxFZ5vRg/h+C87CDOifaFUKtjLv//s+XgacDM6p/FyuLLeZa
e9mx4CPtTK3kt0AyVUbR9GilLlsNDh0r3gnr5QoBFHFOaxvIK1MVmHRXLnf5l2d3
g4Cdt1LBvsbwY6uQIIo5Qf6tMxfhriZSKgNmvWYQlfgCCMJNu98xkZswh/2pFRUf
TpTc4C8zw24HFwrXVuJkTim3Rk3D8P+kRUeY2MDxM2vaQ5Zg2ifyaDX2hFByELjx
u0HfCdsp3eS+hrdNAzKzbff8yI9bCi9NAJipmgVFRg1j8AEHURkkwkh5r1GwcMZ3
uO7M0lyEM3Q6kG+k+wmPrYu+n66K3FPlHBIAPFG3iIjtSWzFKLNiADjup3YVfb7N
0yE9TvLh57eAHoqHsjtjA8LpNt6oCYfALU5PZJ3uEAbCCFditSKbZlrYZ1oggCA2
W2R2kIUtwm74md0hyaxvZVawZlBhEQ4kDkGcpnk/avTYjLzLio1AMLNtd7zt0Eef
qxUrvfp418E/T+vQujwDJolQs6bdfpdRvj1Drz4o9CVipJjSYWKBKT3n7AZPLWHW
mFTDwSObrUkeopXuIJ4ZQreYLBadswtfg2wDlpyYOIlZTEGKOf9tGGd/qpdDJiM5
eZR4lDEMEFrDn/s/ie9oaY72DWtCAG1fFWKQOybiEtL2tLhNxsakJ2kAI65qmrvP
8UE1hV3rwQr4ZKkBf6I6ftVSJnlM5T0X+M0B1PYj8LdyRCPjlMI6IzMHAAam8IFz
mHm/ms6fp3e37Te/Zu0tcS1fuNYJz0gSt2YyridrQhKvRLCygTWtJK6Tf9y/8uLQ
ONMF7gfpkIBIFDV7makkAfGWQWN4Ndb7Dzt1wHL3IKMkxCKPZKaK+BYQu8YPeTXM
YmDICbQcQbNU2o7tOSASZU5Zf13qxi0zWrLIkLRX1LHw4nWoJS6/NXDjv2YPg1Vc
hOeh6GS3zfb5nkg1osjrBB78HBhWE45ATnxPjmjtru8CNSTcWafw6Z8FaoU9hdv6
BgCOb9OL3MYLQvQJtHT2LcenqvKdB0XpjLxHirb39We+oA2XN4F3BFySZl2v0AXd
qDkGtGyKZ/Nt2F1LArUYbkjHUFdAt77GEt7SXMwoodRdmOqMAHd4OSMVL2pM9efR
dbJjxyjPAJNDo+ntVL9HepLbYCw9Mrl1vDeFzFL1qjlpQOBmnxEiRiilqVHH8ZmP
gXNbdb7D/1kjyToH8yVXWIjK80KFw+bKj8wJEREQo/JEv558f3BiJ6IQ+eUr+iV4
2zNMvUoxfas56LgIexBsq/BJTMeeT8M8+aNoESuPezQ3PfaZCRqtPq0g7ZnMUzz3
TtSALd/nlf8ZROiomq3U6j7LQQmC1Mi+FOkbqImAjTpYZvT0pFqnSRDRHT6bmBjU
3GU+IYscvXdrYvGjdLl4tRe5TDpr3pN2YZPKb4DQAGstrNw9Dm5U7SGyz8vSv7EM
mRL6i8Z8dvJ/QMmDB00PtsjTPY7g9hUTJFw9Lbiw1NPumJgJxELTE/3wggL72A/P
q5EBuWclV3yFJngScruOZZLsJnzgvyBFUYASaKTNlzEHCysm0OwbK1J3vpj+GDSi
FBbmF5pNe1IuNUYwhR6XDXRsjaFArMycpJ69JWjhb9KutMNMET2PmchNG9HX34FV
IIjrSMvlR8TlC5gj7u1UPpop2EXmdgKsBX8uH9OoHB9UjK1g5t0osIqN1o7PPghJ
pDQCEYzmYxHnR9xvfPSDtWnjKbOmjvsE1Gm28SeGBUUeMR3dZAZHUKnnb5v2Vg0C
ZZqDNzH+YVVWuQDs/T+XiuSxPqO9/0YG7RCZ3FAZLMAdb4SEe78OlFmMIDNlkGDb
f+iTzRBQlXHSk/O9Dq24UtFtJqigygfV7FUHeTlBpVWqHkpTHsMv8ogcVhKAGgo2
HBzpCvcvHOQkAHSlT2i94IFBdjTYEqqZ3m1edaZeTy4Obl7lu1V/CJkZps80aS+J
grB8uMLGcmA2orsCObF+qIcfvC3MHqFKcC6do9Q6BmrQID0ZjQ6YI60U3l+i2vtr
GAPm+mht48dz3xUAWmp9Jfq9ToQcCJmiFAGnfFc78c1sBBAgmHEdTuuCe1RuqVQq
NKy3eYfqKA6MMbljiXJ3uzt/qV5oMStalgSfYidFMrdpgI1aVijyRhe4CUpCg/tx
GW0WBKywjJEj0izfgAilkg2gKw6YV0QdMK8bFamd1xVA8sJ0kQwZSkciUmT/X6C4
D3F/elUN1IDExMt984BswRPx0Q5wVFT5syXL02qieJRyoSH+EkVq3ntzfTVZBP8s
Vt0V9NhCjC3u+eUAWbShNtcdWGEsn0vFujmz3FT3I1GEghDwcY9xAeZTVKhDbz51
INAykJV/AsFZEFnrjNaUK2Zq7ztUXz07hFAhN7K9cmDXPWBJ5YRjFxzaZcsCbllg
edm7rlLRyZXoTsblI4mzdIN3pmiT8/Ypn88BXQRAV2SFA07geDvjU4qOnnVFt8qa
Ge5x8tyefnj5fRFiNL2DhgZwH2L40Ujabitmtn9Y9XRSXich8/FzT9sBLFI6Aqgn
bjBR8vlqTBnU+xnK9e9ObsKyLztb6Mj6upiOSSrma/HgiSIRW6A2nSaHrX4CbD+Y
V5gG1nAhszeX3JOyTLYg75BsAlH2SUE1weUPxZb9Br1ckjyC3oN9J00URc/MxUWs
9Rt623oPSJZMLobp6ziK/PuLReDhHNgdEsisaedWbj+Aao0CPZzhNpDR7gNitZbI
6lHwr4Y65DzConyxqAq8QpO4naeWzheBfV43QgJehneJDCiR3litvLrJ1vW0UP0i
7bKMc7uYXXyGarJPzh5NnohXaiVZ7sgUxK0/PheqTCFf+4Spk07nwIK2xCpYS7DK
BQwJLBK4yEp3Y+zFWLkXRDCEhnyx9sQG6jy+Ot6muZA/zSz606kcT8Olpn9LhpD/
8d2EQ4WOBOBSqXJX04CCPbBEbVrR2n5dUkML6TxvWTCqTLVSBKQ4azmCCQ4TAlaH
4qHvEVsO6R3XG74A3PAqO+Omwhv4XuhKGIHHRwRI1sH1HOHw6ZTQG4hlzUyeJxjq
4tdtqs+wyM0KkihjnsqDQkiXbNa0xredJ7uHryUDa4P1y+K9o1AVR/aOYSFy4b8x
LY36a7C5wAZpwhUyIJ40hA3NTSSb8731Ie+s8K19Qm08O0s7Rwxqb3jxDgQ/oHvD
Icq22UYpV0dTQXJeb/cnzhF+LEmbD12w3ukS1Ky5JNXXbWcC91/6i48BxfhOFaaA
tDh5Mt7/pPkefTOTLxPWCEkxFCbvuz6XfH8kPZPqIy47mxZQkbMCyTJTKGOtcfzu
GQdUvZIC4DsOQk0JOpaX5fixIKgDTvyx89mokEot2drlkW8cq7NP48KqrcEhHs4d
jfjz9zTonHxaPSZadOTjxWE0HaH/EPUxHHS2hfDlHnwgQqu4YGSCnxywVI2HScYq
OVdMByiRMfWrpYQyY2G/JaDHG1l0llvERsvddHGUBwoaTR/EtMLY0thuxoVOQIIp
ovaCJ5Ct9gIGPG6musBnoeClXJcydYeYb9oddvBEDgRoGtTqW8UtIrhHy4bgZMy5
OECLGBNgOR6dfNSUcm+/iqPwvLy2k7ktNnSmbgYrXFD2qGe38K823ZL93BWqRV3D
BpLxy2bC5u8h+gSgAKomOyjPTsixFDnRKA+t2K5FNxE+K9d8+9BXcy5aXbZR/Syb
HuR/QCzRJ84WrgSfNeWQu8cujTOh/lK1NDuo/zF2NP3Vm3Jmu5XbfCfzv/V48yYP
/9jPxyXCgasrV90gqoH/0NE6QrvT8rduzEfJSCg7pwHHRuKNtjAQIB71J3OV4Hpw
gIXa5F8UOn/6QwvMN1c5Mu6e9ZALvmOmTj3fNVtqAQ6io2gmSuQztATbVG9eCh+j
qfemxSumKTqsNsquuuZSKPYweHy0jnjyqd4LcUsOKLXta0Fs3bpobJgBL73t3qsc
RU2RIIoNiQtMhwMsMaJ4Q9O1vIOJbmeryazHhxEStB0Cy0ELdYU3V7TUY2XfodPM
l2fhnc+LsjukuFfPkbuD1T96RLsKhNBIsTh2yR0LwK+f4ThdDfQetULdZ1GrSfLC
b0wd789tBgQhLX764beHfDYqfpF0+Aa716s6YjNRgunNa+inXAg/oeaJukC+8ij6
mCLhgRXwP1rLAa38SrlgI2vHDkK/unuh15obgzYa52yZdYeSAQA1EONe+UuC74io
idfv+Akg6XCe7Mo5J5FSjTtne97q1RlB5JKYntkUBTIAz9E6oefG9X+bn/lPxtsg
UGSHKLw8p//u6KEavTql7vR6EujzC0CjPTSjF3A/C7aXMlcgZEBIh5/UNZMGx77m
YIIRhy7Ln3h3FTZVKje3IwQnn5Bl+7e74S99tU0An7OBzyKy6bN7Ue/Zx70kXor8
j4+b235QqcUlyMXCDwOYm496jZCl8KlF2yEa5VCZ9aVFV4zN6jTgj2jwOJsp56re
mO84ZBr5jNhJh3dlWjFgQToMODbxFNxOa0eF+es+ZR7394huV6IxgPaXUHohxCoX
6+7swzD18yIDTZWNMEm8Si+5fFYkBEh//uFsgWufuSeFDOQlzp3VQ60v7nqS9Rs6
OhrynJg3WpN7PV+V+ecO9GMqDv8gRgsffnDgyM3frtLOqrR4yPRf2E/AyRQVRKuZ
7vD6iQa2PxjQlbRU7LZrUm6ue/rbsPPjagrSlA7vP4WOgVkQm+h6mBzOAFKNtOG5
Z2zegwHbbUmTWDX5Ve7yOXttOy+pQtIecWzLy5TjbJ+/mpMg3qXELuzlXMQrHMre
TxGCqACl0930vWdDalEv6IXHxsApRwXYjC1zHgjAH3DUW71sRCILVMv1lXxOjWB5
KS1vauHf4Gl6D8xc030l2j/Ynj2did5kJ6nKd4UsZhOHNjFNjQTeum0Lzp8SnNB7
U+i/tnfmIrWu1K/+SjxMNvWtXsMgH5pogPdb8tf7bf1HUwwIB/pinlwL2N8oyMgv
KJZ2Yu0SqZqZ5rUU1ZS8sBXDBKce+qDdqgVdsOOuFjUSPp5GRth8uUl4Yt7NIopT
iFGdmQ7ic0wCX82q+VFj5sBL+pXL0kj1AQiDimbvgtT5KlNZM8rgpzxoeIoKom2c
Snk4252Ff8Wgy4MzN/FEmOORvAV+yISXXGoHRZYZeoJ4JDwCTUck/8+H+i/QKJwi
dLzgGMxR04SPxKLuwfeodm7CN9ZJAS/f32r4F109bFLJwV2g1UaUshSFQTRPgZ+s
KWzq1ZhUI+FadRRSR2JAm2r1riVJKkJDSKh1rrlUVNm/D/Ws35dKLixg7XFfVfVS
88Nl63QXxu+dBxSHLYARQn7HlPBA8rCHeypEcXhVJYc5UvArmwPFrLv1mZOfS4q8
0I65ghzinhw4DGm8h3Z1+Vxt3xpAWanBYj1TNM20qePomY9x3ECpvtmBwcYG2OJx
LeAFLDcax9613a2Prr1qfui6XBHUQNQ53XcSlWvgGasCUPjL4Jhym8zDYeqh9Z6L
sTkcBylvNAVe09TOvMZAWI4QaGNPnwsDa61rjl+j+tVlagw9QxDtNbqYi+FRfVNG
rO/XjJUdN6rXQtxe7Tapdi5UlUU7a03tsnW+yPYBcRJpNy6w4mGN3qyWw0EbajmU
5JxDG4s4SgC3OntV7DE3HTsRULe2VgXLWzhjCBMYAvDLo8VmQgsOp43oYyyPEkk0
uxcx2FKSWVSlV/7xUHrKg5rf4O72nCjq/4U1xoE4bOzn6fw5LOhLRGtgyOQ4idey
zrlYi+e9dcQfw2LpNA5mJm38CMkBoWGCg4bXi9rr6nq+CsJzXIXnEcVD4afUNj74
mwYUMDBvQ3hRJfFzs/ljonLDfED8Z0C3cO69j48TxWqFdydIfpVT3/2exF8I8N3o
JoKPXYyAtpk9G0chSpXfZWiFX0qTSyOlRr+bTrR6LczNkHgUtEpA5q/PZ7QRbfvF
90fdQMzKYVODPSGyq/kdXVLfau8aC8KqlZkkJfhxXD9ixEmO7yLekSSC9g/r5hQq
Dilm5W2+7tXVSA7nTGfpSrTDbl381kz3zhwGe1Wk+K8IHvN7GXzaHqeEA42hCBkR
fvIBWLgUlFo+KGXg1sYAvpiecM1LNDAbQML7cyPbNKmmon4vozDc9zkvXf3owEfH
aT3rZMjnEcnUvxdNw1ZGb8Km07LHAcrSEHiqYQN6I+j9l936lXwiUlxpsEh+h3zV
Xv7mcHL4Ya8rJzHMC98nB1CfJtS1fZdmovMY+olPjbwXPHFcXwx2dqgaxJ4AJ/vp
bozDf8r2cZiUNGKeMgWkzfzeWqSuZLe5nDxUKIN9pOmHM6cN9Q7idwqRgy5I1wtl
q3b0LUrfqNdF/qlPvFEOiod0coLOiYu+0+crmxr5BCaEGgc9G4iPXshrgAtXFUg9
cu5V4FEd2pRtJiNSmlRGro+Bo1I40r/qcTg14g7c7AvFfRRN3Max3JlQ9xIq0XBm
DMKkFQyb/A2FuUoG+70O7tYdfU53nV2PUKW0pOKRR+pi8rpKuf2pykRIzTMY6B3T
N3yZ/1P4Djr5vC9M3n1CWEdvbmMJazXxJQuMzJPIuPLVlEnGsNxzKfIzlUFrHPEl
h1A+skLcAXHIjQwRzqIrDwF+Vjv766AhpRdajiaJhbW2qVxSV743n15GU8k7bP4b
188RQOcrPfKtGnDwk7+tWLMpGrLQ+o397gyNPhprO6U4fP1FtA81C/cw1bjJYMG0
OPaTCnmwWP3mMTZmdQvnZNmaWxI+mSr0MKs9w5YE5OypguhrQCJmRPJ2OaZOUrmE
iQXhXzfknYcLOzEKlOARDugNt7n4pQ1ks3ttp6v7neBhQNz0M/YtGgKDiStfR+rS
37XL29gzqZRBdr2IkUhBnMOdC205GfEzPUc4zQFP5WFr1YnFk78sqEOck+vAEFUD
w7qlJtxQm1blRRhZqo/OWHCo5HjyDt+DpO8yQTaWpwima5pfjXxWu+zXTmPGNjXJ
QmvpLerWSAFzLtm9tc61eNBIdCSIRpNqSx7r1LWMqTyssh1fW01g2WEFhwCobxXv
4o/6RgUHL67Zo+BY5JXzHMIe6JhWZlgF/odGxXQeuAl0ygNm8wpvPgZe2hviPEuo
Jiu9QxumsSa+j4mwdoOq9i/t0TMug8sIE7MPQN2okI855dx22fZXH5fZLGiEJMsR
RvAADxpxcdPQx6zw3MJWEEMmycrSLijrISqkTzLBNIraI5JkLGud+/KdvMrv2EYx
GMVVBSJPeJYTFJO0SJIMvfX7K+LO4ytE1HaBzcMrq3gxzt8rzFdroFkJFRmXU/fb
Bh7OE3oUJ9R9XoIVsglgjqvIQRt5W8OIU6JhnCjreTNEalHdm4wxruZKpqHOnI2F
GlSXMVvfuaQhkgJsWt38jH5xgE2VkhPcNg6yWWXkx/jbv2dicDL12ySUlTPv64t9
yVWOobPXhRI3d2RrpGNxxHiMkRPyIItbElpkBpoG6GOPa2n6zep3stW1J7YPH/6S
mXe1RTJAQkcbIh1/zTpR8F2qnygMYkZ2vgHQpGhtuEvHbPzjDhwXVMaXFQ/khXdM
FPXEHk8wLlLWlIQgKyveb9U7rU+sppDXI5+YXIdkgkp8BeXl+Oty+GpklXppfuKh
LyWGboW9T7Dog0KdidgX4u8xNau0rAaeBaA0RT4G7ZV5tDb2JtGKLMN0r98WfJmm
F58OORBsTawyDpNPVx4ZgFKZlCoUSuCKgcvl4kENWK4s4yGjZC+jzeaB1nNxrV67
cv+JJdhLnIYKe4erA25pf3WWiK0luYJWR8YAcDUStgdnzQtti1g7e4FJeQg4vfqi
73umYHvvI1CDSoUhV8x3M0PDP31OUC+tQDmxud4iLBJQ/kRX3u2TAcnM7EGgZNG8
TBPbKDHeNU5ugtAeknQAZVIS1kESNF1GFDcbJsfRUz/ql2vlrAGLITTsUJ3Cf5Tz
UQBms8gu29L4tOh243bH92u7U/2iGdlGn8Xcfwt2eh4WPJxiJQMQrNJ7JkRiEbn0
O585LDWvIb4pBv/Se/BH3fHQeuj8k+YucEFZn3VxUn5+wrt/LhE37T2UKiIv6Stf
i/YCZoCNccJPISCmOjjVMjBgOEzBJS7Mtt3av7MxqkDTp2EzEK7i24sLclYKjLz4
noohr8YV+j8lcQda05mPHm5OZkoNvxQNyhJts98mowBKnir1rMOm6Mxo/bfJ7PPp
e3zUv+Sc6+Yf7pDq73QA4/9QwE8QetUiQDQFFXe0HX48R1mTb3Gx6j6U7OpWCLAN
qngrT0ijF8IRd8jBQF4cUhJoqWz672Tn+OZPSOHayTm2YxLYm/O/iZpr8TTzPwMK
Mow1Gp9C10ue3A7knEExhVc3gn+aNiwE+/g78QvTaRoMpOE5WmcPkmCkelWI9qRq
NohWEYlrTbATwQo641w58m9VK0RARPl9BzozoKqkVJiBqxaZF4IBWgSVlPuSwPye
tEIM+8liDVq/uZ4YtIDuX5rczUi4dljC3qvfEBCAUVsj01rOoTStu/5ePSr/FNBj
7SqTY/SXuX80Bj1uMrdY8tbFqmLys8+XR3kDJOozBWY1X/hU9IB/nIbbbLPF+8Cv
ZbdPRzW+VzwGd5xA96o8jWTstRCyvrDT9v891fKZRWPKZvfNdsnECGE1ZGN/7xJR
sIUfEFHUhSALQwUnA6l1/gZDUzHUNRQC8WjWQceZkO4Wys6538dgAKFfkUxqmVQx
k/7lfL90fRI57MqC9ELUkm91gaLcY8LdHbY8eS4gBSa4aMdYCbn8qozIxEpPVfh1
Vqm8voCt/Oip34vmv+A5fz/qYEjLK7riI/Zh79TRnSTFN43bY17PFS1jx/Mda11F
lvHpE7PaL71GMgozPi5CYjB04rkaS6TA4tXYAwlPYGvjBJisZx376w0rvOjhIlYb
ZZXkAPwxFBhUcYCjBvX5+lwlKs/Qj3tMHZIShxvCmD0owkLpLaZFY7TbGFdXiLpw
1E33LXwfzeMeoDitczNEk5X/J6XldZaFghYitYQzIJykYHeBlyzwpx2Xzfvnxdau
aWMQfAJBJDqgH05X9b5fKAZgth/1jpfklkF42tHTdbRPmSY/9+S2fim8NShmJVRh
2kr7T/yY5ZeAG2lOdM3hOWm0BQmWT1TSYAsw8bjV1job0YE7dac/wgpNEFqujS7C
mdHqr0RDwLJGFB9ShuAvML75DzwVfjVmjNtqNx9s2pOjgkb9ie+cUlreEQu44K43
6ONI45ZdHZYTPeQVWx099EusTowQY3fFAerwm1/lSoSa1pGYDK4Az+9fjLViC2DY
62JhdNURkXeAy2A9z/Q19le71cjmQyRpIE+xF0KBmnwzHNk89CvNr8/33cdNjY+u
ThV6dj7FwTyqmSwI+xtHfbXDKfOi+kvIdJQKu1QauicbXpRSGKLKi6uulpoJHDMy
O9fy0Pt00CScGxlfPaxjXJFIi1tnM35dDcc+gNz9ieXu6yOpSvzy2vdBiomRraMR
Ohr91FEmO1iL8UPEjgplFjxV0rgvdJ1IYJpkJZ3o7kxFmGwmKIN0+XxEgBZUCpjO
Gy/KxeYPdlc/eK4ckmrWQy7d0/9dvQ3bV0uL/n4M7Jyu7ylRzXo0b+NwTAJ4APR9
Ka/ew34HRyi8XjM5rwSbpKZn/jePhCF02nHH5na9wkL0oAYtwfktf/T7NT1B69Q6
lHd47ZK5duVyRcPSBbvlRT4csG/ZqkQq0zRJ1yg3ic4yfqENnMab4l25aeZwajAS
6LNrVPmNb762GX2kvE5jkbbLRJIPHIbWT36sZmbtuNAtHr3idrBBEYVqyWVNllGI
jur6uuRDN5JFtAqtQ0bqCgVaTMV2LTdVXszXl/ZVTqfFjRnFDkK305XtNJlhuFPj
lcFNpxKp9JiXfiBMc4MyDMCSvyncgbEKxGGBSXTRDsIlo87ifUQvURvYVLQmgVue
nhf7ab3ZrPzGkuVQYh0hXYWk1dJMg4WTUx2mWjl5nYMz99CiEU1d1GUMDsfyLZmT
yeaVvObskP9M9g6RZQNJfsFEugGtKxS7gvO9faWxJJ/SH7yigfWJD+udzZTDjaW8
HFGqr7q9/uOd9NFZobvVNrZdFDYrlEEwlq4mL6i9vrt8gkmK3L8vV0OSAPKJwPh8
JC0gEF8HO80TEYP7nWFOQZT44vMsGFn0+UFvFMxoJ/vE1MiUVgqUQN5uQMWl8Jo0
Z5vakJ7kt91cDSqLgEQeN8L2oL7KM6upq+elAKVIvYRzuLqlpcMPImATBYTLHFOj
goxmXoeUZ7kfPUxhkhynF+DolfrypQ1aQ70TDBO1hIA2v1/+68jy8uQhWM3gj1bK
ikUuz+5GSz68IdiBSnOMU3VjwvymgFw4s6GIJG6d2Q0idrNlW9N0XsEQbeNxrCHf
sz3DObeEQxMsb1OhNH95XFH37y1dmmBvuBelsL+WGe6hUK98MbZ6bf90MilRZVMC
PaKtToPDURVaEuOLj2LNOIsq6rvUqS4cidpZ2F9AycDbEHT0BbUpvu7hctRfymuV
tt5D3hGHvdrG2PqWpP7113o8hwz0zoYRu5b4DFmvM9cihjV97L5B8xrRva9z2WkB
PjgGTg6UqFnaAnSOWz/R9KnJxFUxqTeblcVRB3zR1rhunVSzr+E6PWOCSVjE0QvC
Y1lPd+UpLiIx9xdj/VMrwXb7j2ANIMU1vA8EiRBDSAo8BMoYhdKeBNu4UBqRZYmB
W6C5/aNplY36rBeAboSibimXDgZF/nxjA7pbx2tDswlGpzWbjz577/nEqi/H5EY2
JGaZM2j+8aR57URSgV3301q86+ddo14tGzHs2gudyIUPxw8bM8F5sdxT8Bj6MOJw
smWnOVo/tnFsK7mIWrHHMf2GuuydUra6Ai5fvWY94IsXQ2y5fZ2eXQbShI2HysHn
f4SE5FNwvP/0N2cvERIASjdozV4LTL5sjKnF2YizwrwtXIyLAGdUMCz6o0OmaaiU
rrJlFaQFwj4rFuOz/SWESX+6iktx8XUUVnz3rKMAVSR7G+gvhBTynmJZv2tfvLd3
1D2qTsjBtUCoGIeXXcQusfuB55qck/ga+F24AQ2qzuQ42P/9G1HrHiV6T3sQGvNV
wYjRwI81rn201FUCGDdQuwip08V4a3FVefccnoLfU1ErzqISDWH++GgsSaF3cq1h
pyeOIXh3ekrkQ6QD+QuTmK8gCACbpoqjWtqjYgVgjxQBtYkLv0u4dTlsXZyJngDf
qqS+ECNsQd2Sifddhu/BuDbtZAeCYENuwCJoPn1WNi/zFJIE7g73UKEEGIfRNact
0VXpN7lRfIeHDLKZEPTPwwQnXDhyG7Dtdwhnn3Q3XGieswfl81xhkZC244VS0jKU
0+13eEhcqgoaJdtc5Wbq0tkSrlTIZTQWFlPdPmAcYq/bKev6iLs8/1FReMU67bBu
WkS8wwY/QPodGmSQsT/RGBjUtkutYYn1BZVE1+LP2B8HBz5eetzWOtwpG6ijq4T8
h/McSUS62Mjl9Hf8OBt/iL0hArlBUrASs5oXCpwQH/SuoD6sHEDHo1l9Pyy2Yted
T8aeKwRFnFRCi2lZiv/wFVGZyH0NdOaN6BpnE7txi86ePjnSjfY3ACaB9YUxQjFm
uzGeNf3Ax4oMNegKE33ZOERNw1lvprOO+J+gaRq1z1Xd9r3w/EYePlb76H0JTRlU
yqJBdZBBsH5zgiSsHXnbFER7MZSuVmJOjRDseQvIDBQIqQ9EtYR0qltkCAl5cX52
Ckx9EpImVZbkFpl0Rtm5u1wRx6TIOCye3Fljg4a5RpeALOkdK9BJm47M64hjUD0N
yVrN0HAalYga97YeYvwDwwLCMdF0O4UynyjvnTV35s6yidAah2YS+BEfyfbjshKL
p5wSkmENozcAhAcN+Hqml94drW65PX2Ely/TBs18owTcacv+ARLLXQnn72X3HqxZ
4ET9m3IiPCvYBrbsrQL/5laiGlVHA6cA5Fy32q5+8P/5CoZyPw521d6tgVJ+2lVY
t29XDB2Zci6GLST8QNwIkNN+3QDeOFMRXYs2hJQXcwOCvd1e70VjXfvPjjM6b+s7
lvw0igqFXKUfBiUVvIpS9gnUZHwINZ3fteTpb6hrpfgYKlY3/x1/rlmrVca6jpIP
C9LV0Prjfff0c4Kkp+ED4rwbFEMqlg2wfKsINwB5/WFIb+9ebi8LhLWyPIO1SVmV
ceZfBHcR3nqNqmc2hOpKILN3BNxc0f5GHjoP+1EjViv/N/8+b7JYWrB98XBp788O
7Ap8dRoutPIrE2ZrL11orQ/JMF9fd3x8Re96U8iY6p8VTnyepziOUSmu2RQ8yJ2n
yZsWs3sX+IZMHnHgmFk0vhxEFC3Qgaf0kiAcqtLk7/DGWbWjZyjgHkdH/4HQsCa7
xBAubDm7e2cNlfqGvQchM+E3jXPyXlWzoJCds4jFIDEdf1oGlkjqXESdMS5bsyE/
GMqRc8ODL6JXWECeOPZ9Z5U51QD4OrLMfsYzdPSuKdjzCLBUWu7W842PvQiPPmJ8
VOyyn3QM2+3qHX/ul9bFStS6sEmfn2VSd5ncml5In73j8on62mAqhP9m9QjMQAP1
wwk9yj4PheK2HyfUuMDizTj/v3ceNo0CbXVgr9nrSb99qaPdiVdTBLhbmHNPFlO3
ZDza6xiKGIpSeXF77MACfQCpudhvXq19LTqkjVsPHaypXnRVh2E6m0oReVTLmeQu
UUs4SysGzugsI/SWFy+amip2pkGmh235OZJ4jfKZTyoUz7hJh90X5hBSaVo8mcTC
/VwYOnxllh1gDAxXAUshlqypDE8eS4158dzoeBVv4QWg4oSYIP/P2KcX6+TDTY9F
voNn7fFHs3PqX5hqemJtyKUvuZI5DY/IT4wjLvn/L/ARk/2kkvqMc8RwwLepVADp
5sYL6YA6s89P1Oyen2HeD5DU2M6jtYihcfMUSVEBF4B/Zcl5/BDuFtPznwACqy1T
MV4QzGFuibhdYwaBWnupyh3nFQHhr92OZp8AR/Oy8VL42w+hXOra6EBVwIxZKFGl
TVpqT5+2UfSvrYyFyYjyAhqueSiPMy2VgGDHYNXcMR/b7yf9IDMapD0tOqaW5Pke
eIbjAZtr1Okx08fK7NAwgRqVLtmajIOZdzbfIs9A3iTIFcf9/cumOCGWxdZU08qE
uYjOXbIDVFgaQXHXWHE9QsAxWPA0/OKdC/DSA7nOXBescO4z2Faf7kriirkIJBBS
Ayf5vPA3kbnF8leByxOf7EdkLWjmtb4wAWusH0V2NakGFOZXpBehTT3pFIt8ySjj
k5iBqWKcMrCO2DA6SAb0uWts7sVKM1ji3yl6DIZhVg5ApBdhwyFD568aDphnXPzI
ocTr9ChrtwczrJsn9akyZvPVPzzDpXrIasvn0mPQGHILgJ7VekOrvDPGgCMztw18
FWAY4MQgXBCVN6zTl+vs1gPQaO32KGAJrGFejlRBrdN3cPhOTKeP/RBJug1wBXYC
wvyIXvEiE1BWwrogRvtpodn6vmfngaCBpht3plQUje7RpE8Qqvvp0aHWiYVfyGRi
R+SwZKis3TovQJjzApHA7/xRmLOBg/XMq/xuPEXgjEe9peObOggZcjPeWa9p8FGq
bkApaWWivGoIOwu9WzEVvUyi4E7Ui3dEQE4G4ze4GAec2day9Sg9h8pS8SbH3AlK
jydLjhw4LVXDuLSNNwDsdqmNSnsz+bSzoAXReZnAvCblnquBLbKpvHCUs6iVUEu5
wRMcpNOhnN7hjUoxxpva9rQZ5eFtSohyioDpAc7mBtWQ1YxkxGgejjLPUADP4JZS
BlsPhbyIPCGR0q8s2Zi/T62EhXFrGb6OaMZLYquNYrqc1Gd4dfEZOc+Q808FQf3/
eGuwuVv+FbQcgwfAIyWMGq9watO5UCf8ABcUdCC9XZGQJi2MnyUm+j6kumNmq+j9
KjKWL2NirrTtMI3TRSun86FjRge/h+fY9LCK+6NP7tXFXplqJh4iOzE4tWa2VGOm
YboNgR8L5RCfnB3GCSh0LSolHqeyohLIBw/IXRHIn3kLugECOkTBwLSs441x9RTm
sZwKFnSOXALoZcE34kPeBVfgzvlM8/+qLCU6toKCe3S+RlvD7DB3KeFw24pZLTfc
oDF1o/fYGb3Pe8xN+brEvDBIBNpKZt8UWlLDVhdpvADU+ABZwbn2fNtvfAu3s23s
mJozC/HOkmGKf6vSr3GBrRr6HejpzPlZIXpXOMAURTLwp8T6wtQpj3eq14tLdCYB
wB1BJK3ZFrSMAm1SVek6GjMcInXr27zmWemKI3CFILaV2pMWs3EDFZrCsG56d+Nj
TDQM3L2X3P9eAndKPmIKClIFgbz1YrE+UJCIHEa/SBui8WVnS4XBAKC0AZmTlwaZ
iViU5y46o+/ESaD+/5YynG45BwdqlOXXXxurhwobRzCNvzvwZUy+msXdG4TDGuj0
dStRr4aOY/8uP1mTNob17Zif453qD971o/qQ6s11QzQWiFxUgIoNHM1POmx5h5jn
mZwB6dHdUovk33J7y2HdVWDYQZc4A+vBrG65mraF5stvRzJYJqd8xI4hoXvvL7NA
D1VkxQBNJbt4LdXYF9qmIp0YnmhaRc7m5ofLjFomJhuI4BDpUX89waBp9cf9aY1L
iAKUyVLLU5r1VqAEPuoZMZa7d06VPBxtjQgPnOZKcjIowAIdEStjASvgee1D767S
kgnL9WA1eiv8qk/VDtgAQJm+etwMlbkOjvDhQmVO4V34Qxhr48A8vdfW1ZJ8rfD1
JZT3vBfz6JR5WdxgFiumKN9QgQTecoS0bd1SB9vQRVwpHm2jY5qZBpJJrooHKdI9
XUd38N2dDzTTVHBvlbwl705hzjQtWA72iDv61ZE1OEjVUFaKHpz66h38BTFDrJq1
jq9fnWZzhpGg0Nh9yFdCpLD3Ie0BIf+TdV8Wf3x5fTLcB+H4pt1JpEf3EuOCurFi
TyMhegrytEEXa3ot7cD0SU3rZ/2yLzJYHB6zUbEKTrbBAsZxwsnwEB4Kiwf923/Z
+FL9J9fSUMQf5NJMDwrr9gpVrIAUEU0b1yRVFXGHZj3YfSo4D3jHcXN2djLEbmAC
f9L7cm5k/e3981ZR6/QpKHylMOoE8MuSk+Lft0rXqnx5SgTirKF/C4MnSE7TKqRH
vEk3tO4wn9Btf0VPdnWGvveIWOnmrU3iJDxEvG0avrKU5DqAzW1u9kBRi1czExcI
fva2ng3sJFopkub6XMHooPmj0Uwj8H3inYUJJSoOuWCliAyfsx5APnnJjBIXsHUq
5MbSIK7VfpIhrnBGY4oCBXgBXIoa6nupDTnH3pve40iVj1suiD4PHlMMjrDVjyRT
h56dGRDcQF++EC6hUfzNkFCogY8LbLKgQTgoOyQHROXlGpyQAWmMT6g8TjGh5xNW
EzhFsyGSqVZDpSGTRo52fTMmj1pidqd7xASP423Ma9lUrlYWmQzvmtDmzWBhJ9T1
kEIf7qkRB38z3lS2BpFnx8J884lt14GLqbG6QvTZoJfily1Su+BgeJi7MkZLQRkO
XqbeUvWTOASLlh/U8ut6rmBHieTWapqlh+wrLWzDHH0XqmswKQgnxl1yIkCcahDb
JC6bAv8hgHUS8pwOm+SxJPB8Uvikj2d6ktCCdT7p+l4EnChTFptirAbZ4ZPguEqi
DJSyNfG6wvuF/0bqP7KRrykcTdBGQ5CnAd7IapTZ1nDM5J/PR1Zm0uyI2RdbXMcn
zn23KRI2rxHhFfbDEC3jFVAtrCmjcwJgyndDtktUXWk3krhXtzZMmOemSCHhprIu
ilsbcmhHR0W6DL78gev6qQeosFIojod5j38m1eH4fR7t86Dpo46SsFPnnrU1H4Y2
iqp+Lax+LR0pc3gZhctGBhAYShYJjlNsb6Kv+BxM1geeTqowe4F66e7IahAaJWRp
fgJ+fxGq39iyyc7DGezu09fglJWh6cZGPesuI6R69Tu/+uyJXgknBRzypb7H5aTR
EO5miBf8TX5qrIX2+NJD/KrIooigDjOMnGdi8RdGjol7yqvAjgkrSeBuOLDEg/YJ
/KI7FkSVKuztwqhS/PqWOzZDEtgYfOrtVcqCFH3/Vm9WDl0q4dQ0QO90J2c4x6pX
sVHW+drgcBVnxEVM/V3cwKzDvscSo+UtFfLvR4FQ2ln9nxi6bQQOeuYdvi2KEkUM
VSqIkUV6qCC7a7KtmDxySip2sksq2aEPPVHJFLx9Aqo3n1RVwV0Mb92eCKSRL1DG
5NghlnsUu0xKFPyEAVgO/tr3RNQufFZ8flFUiP/yxYxjpEtXERawTM7/O9pb9jEN
2J+w1oLW6eA2xggnEXpt0fcGVYiJn38dZx7Ay2DnkTyEkjGJF0TToRlGV+DzolJu
yEOMIlskfl+jnlLA/xoc4EZhxOHnGDsKOOA3k7gNc8hIad2H+6gc3HFnPjAj1JQ6
uXBMCc4qGP0MyQcPzeQ9UExWaYCi3QnYlVn0MylIGFzfI+H+QQuKM1LhqjocB+AV
FD6fJG8lQQECSehG3KiDCAqfIEaMveAIKsoIvX/PMtwhjbCoMOIucQLLHRIKWL2a
uW6k7BL+57dV5IhGkj5a4pew/serjptkiiTJZHmAP1P7ES3THYxdroA4Sxxpq8Ur
+HAEOq7qlSg182OosH1ZiBFs7j5OU4gyrUPKH4YdkqiwRc6XVQuyu+NqvZNSWol+
B3VzP3FiGHg5a8C300N4gLROzQp2SNADVfdF2X/zeAzkbRCdks/QxJrHC/LLL0Y+
B0x/geVOFCh893LQNNRIiGw3Qk2hHKMu8piwJCy1vmIbngIK3WTstjlH7nWKkzmy
HVKykZjqQj7kCjukfjZb5narAIY4DpQ4x1hNIZyjdSIbIdlAU2vGRMo01PgfpBfE
zPDDLGURERtiY/ZbF0ahsImot98lgOTtFqNYwciCjGPRjz9X3m2guPnVXzkuUdJa
vE2yoDK+1v87Hy5+4aqVd9Nz7AtHRTU38Wf4gHO6Et6VjmUm26+JA0WNTuEJQRQF
qstgU3r8Z3zYRqM6t3ti1cD+ryOklEXORQTqm9WWIx7eD5hhZeXiosWKCfkpLBNY
CpnLpo1XXIAbQR+Tje+KrSpoVECVT0pvCakH8N0bwTj3QQnP8mh7ERwCI8n9ZC1o
Mu7qtLAlzv5tmZIr+zqioMPDvGyuo+OiwYHw/EZ9OEZ8Ecri9uH8BpdAtnbinYkE
2sh466Zpqn3qDebCf2N6Qfeb6v78B03UP/Qe6RGqEPSv6xIonFm2r20MBcW95EoD
obiDc/Ke0SDGOgSZIpF2ZOWBxJ9l+FD2MeEDMJG1e4+hdyyVdelITNHq7/O6WuME
ArsN7zQCyOV1waw3JPaH30AS0YpENEpmqNgZ4epDmfJ7mCSGiDsresJ0rH8blQft
U30CyfNa8Fza2fYb3XU1llxFUracwQ7cxYbkxy3Pmy89MMB/ZnkxNpyqrU8hLk/1
uG0EUHOO2d5JHvjPhAD8qV8PJtDJzkRQ3p/cUhsTKFvMdjZbBnFK0BS6FRl/LRVu
rH3ue6TzAQF5szKzFnI/C4pmxEuWd/4zlXzaJZQfetLAaFfyISD+XcflRpU7/WdR
jQB7ev+svEkGRbaF8rv0moXlnh+kbjeDyFOr3PadCr2V2pULbdVyfjU9gu8/SYwH
5Chs13kn2yCIVji6ooiY01q/nuChnkUk7dPxk8nc34FxS1xZ0K2HiGN+akgUkrEX
gM7NCCbzRRPfIRDwke5SaXqR6Cd+G7+gMo2GpYbkzzJODYRn/BqnL7buP0CiSpfx
riK1bPATdVsqH2UmD7dkbk8Ow4wdl1Apu11d/3yqhUCFooYlivYi/DcivZxwQpFp
OrejSvkHAZ48aNQLz4kzpAZ4lZmTvl1/2gEqF+N5Qh/IfFKJBwTPpPA4dcjrdvyi
ajgy9WRyPdlmqpbAtEiLdlCUPbnm6HcXnQUvv2RW+v2tTmoPrq2+XjzAyvhDGm3z
lJUDj7BljRgWVpWQV1pgmx0Wjg6ytn5NpU6dJ9qOoU0J0dFHJFscOG3vDBX1KLTl
9KEgnZmvsTBh9QgIBgAmudot0tAs93e6GTneyxqwNfeqBOt+DQ7roB0o84n3xAjl
9XZSgHGW2TVJ7Wa9qUa2bsG3s81i57oVGHlvJiZQ4EVPjgE3l8lNbzKqRz4QNaPw
397wFIostlfkG8ZtZWy5a/FHx5X831Tz/4frUR5STfJ7vzFIE23eOtPJo2PauhpY
0AW1IRwcs3qpFB2isJLCTMp7Tisd0saOSGRJHCkVVOZ6hLAXzyY8eZA2WUl3ri/k
D32a6ClCCEQfhteHCtJIy+Vb0BgaHGDF6hXms3l3IowPsoBxNVO1F7GlJSw+3MVT
UyxYq+BoOKuQBsLQP+gJM34NCKBXTpWrgokzP/PjvgNLpc10BFIOKgvY4nqmLMB2
evDy3ZdRN9PDZxjWPnuALiu8QGiI50kFn8NFQ35ABh61URSMFtjub7PdyMbTM2Gr
M5yTuW82WZz6dWaA50Bm6YIY9rchyOfPwjNUTj6L6W7spKaXeWQUYb1wf3hk5mFE
iPfSCT9NJwkehq9l0spytgFMXZba07E9nKC3qqy4qkzDLG2mm9Weu2f/k9ZJE2vw
oNi8I/avrOUdYRCuWqXZ+h8IWSEzVDzyfXyFii/1kJm9j1QdUlrwj1I3ZbwJwDvA
z/7es3g3s+OCnn/XtzPwVkfi2nN+nxweA+VNjfpSBb6H+mLmaMkfz1jeJmh1b+A9
w+H2xgf9CORcJOtp7rU/tl/d3l01FBnHwvypToMKxvDxE31q3JNpYPryboFs2Qkd
kTHIZSNeOFjpS2SP5bgl6k7Ed6Cb8codKOmKSL/UyH/53I5SMapUFw79WZNBLIWh
VP39SJDk318I0nk4SlW6fhb4MJ5dp9ILZs2c/RIKPT5+jQuoHJcak4Ak2eCfa+56
qb3kM1IJ6GUaTXHgi8RF5OoJXhAgNKZtKaeVVlnZQxrQmuGjdlCYiGDvjiFdwlye
PFpEDXK0iDIomqTaEZoz9UIUioIEzJcvmHqjJI9FhWd2dEJlSb1cEqjGVi3vF3V7
JagTzpwzWKSY1VM1WbGN1Z2znzg9cL9czPkVSj+Wy6GxJTAbkD9VqUIGEIGXY88D
b56JTDvOWciGcubWSgDkrFlteDAoHsAViVWg77ewdAA2g6VtwY0pEN7a8JtrxC7r
rUiGZNJqgjbqyeuqnFRBIEDu1e8zUSywA3xqeoy8n7NtnAYJUfEMlqd8Ve5nfNOF
ZA316V7xf36trrwgFuBRq5zcvLFksZkEWJDeEBd7bCURyfrvya6MOTCPwd2B5qCb
oUeQR3iOl6eOInkHiAG1ventvMFJzPY6MjWxPaCRxx0brus6h86nwoPAsuxYdIn9
0TJcvo1+DzRSni58plbKnZsj++jWEabs1AsQrinmBy9YTYGMith+uGNyg3zoYr3S
zdPFh706J2RZWse2wgd+O0f9Z6wy5h7fNcZU7dOuFgDTgBRvuHEx7mdlu9Q2byRv
3bJI3vG3PvHsULPD3vD4TEugVy1/l68dGvgkWnXZA4nm8CPrPRBtullc7his4As5
mBKugE6K5r74C43h/MfJGhTOnuD1uwc8e1shOH9we1/MTfwSPHjXEUKNTzNCvpjY
p2/0V+Ddou40Zuk84ue2OB+528m9tK2xbvGmeul+OOlNSEZQBOqNyDDgdHQ8u1w2
GPY07K4cthUO3OxNyNp7ih8NGxX6vA6yWbXd8Qrx8kq5jnExUPpKinfUtUErFzHW
BPQw/CegzDniyd2YliIjk4esHRT+4sdmlSA5lNu+GUgkcIRLiiE6kduOMynixtzr
xyOWtDuNdawWEp8PUn1OIV/I8CTTMOMldr9s5rUGYDJCTW4CMlmNHR8wxABHoeRs
Fj/7DaX2/ZpfkFZ7pd1SsFbEJJFwnlnhBPZtvxhMWgalEpGyY2CF1ES7Ll+0Obob
ugQ4LnFckvNnVWM1xwlM06LrxUxysOyddw4pfGF1Nl5j0XcPA6h5kFNsbooEJAln
pp5UUPLotzFTTuNywbegMo826QHGTDrQbBKaRoCVOU5i1YtWLJa+SMvWgKdgWde2
lwZ2Gt2i6ctrPgOvFkB5dwtOx8AGpQtMYUlV7sZki5Yg4CPKywtVANb5SmEv5c84
7tNlEILG3iNq5BgJ1hXHpKRL2FwkAQJJ3j9XfAvpg8DMM1LlzkfUfqYcWfnL1eFy
tTgJzpklYam/hMDVKwjrNBce6Wo7ccZZrltzd2kps79JFeKzx8oboh2rFwRHOSFT
gLqsIw7TwZkPEXQPBsJs/m3hXkNs62hiBOHFrKtUX0NY5P7ZCbUTrkoCU07gOYtg
MW55ejAcAILjFyib2rEjyND3Q628NK1FXScPmeO4/Dddwz3XtKiTjEoviyMC6g7g
plWenIl9nnQOaQGmgeYAUnmObb6bTtPMddwoC+td0th0NZ6fQcSG3CIYxb3vAB+3
Rq0xc+ZdI269PEmsyZkb8AfXrFS2wL2XcARpaLZM1qqv0mSzzTJkFbHir7ULZztZ
oE4OlYa4ctKp96/CA6nIHTP/6YQFBmAQPuOUqzngHc/J1RmA032Q53iYN2w0dur2
T2rZUf4oOg45LzSDgAzQHr73Svj0HAZA3gVVVT7WEsj3SaTyiqb8SlFWnnbV+vO0
SXTjFvOd65P6/fW8t6Rq+fHamni302vMmkdLvqm+Fe+bPmI6HFLfVUTkchzVm3JZ
2xLr6fqnTxBX1j7P9bmvHT/WiCJEDKrKnqHKUv4nL80lCFAqWVCXVnS2J+wr+UKU
CQCSpxMZvFLoE3qVKs8BVL2EqGqN2+VZtYuIEo4rCIMEcbLzxSdOYYbvBiljintg
0V5bDJw0Gk/n4VasIa+CRiwDU/r+BgHqmFUwS7crRqkQw4oWbChzgiOF5xV456in
6OL+XD1CZrXo7LJ1DpMjn//Mb6x3HdbEeYBd7FDC8x/hT6Pz3QCb7+cJPnXYnFSy
O9kVr/TNWzkcfkvZka/lL4kT+xDfe0o1/VQ+NdiQkLrOPqGqN3ixPunZKS/VDIiZ
j1VrZvEmM1/0iBuEj8p58rYm1IbyyQz6WrZlqbz4stEaO5WigmiyfXxCk8W0FnNi
GGTFoDVNVACGVShdUcK614IZLIMyOVpJ1jkj1S8evW39v6YBE2xdbqmGG7SfS/l6
SjDs3x9G3xVIs9J2KvvpnupTQQT+B6Z+q+2NefZztnC8djzrwuXv6c3JKtbvnMJH
tp43tpbA9Fl5hj7V4jzfp1SirNnTNRl9orf6m8alCYrhFWl1RLyG3c/62kzX6t0i
O0vszFJVei54rXQYEhmj6MkIgkWYsuzSaRF18c7QWtrHvKC+AG+KvdNnKIxhwISV
ghVvVLWQoQGyuTAYjqNxsPt0oDkjdRwmLbDlloB0bkxmdCB+eTtpDrJjTVC+D2lP
uvKGT28OIH0Fvk52IjgxfwqO+hjsqLuWohMQ5pVkb5JDfk6zOSe7FryS05ZReP+H
MCBpuQdDg0muyTaavNFK5nJDVX2aHUi8eTAPZnnOu2DQNGeSLAAJqouqdR1BALAn
RwMPAwOBpcga8DGDTRRvLZoW5UggOKFl7mrhUrzFgpijiyn1mgxd3ZckYU0J28z8
h+dhUl2+Ghnx1eOoCwO79japdkA/iw853FJSIizWxkhiE/bPUw8RWE+DfoQSNEHg
S1XYVPLguYT7agRbOFBb4QyyPbbS1PalIqWtIasrI5lkEQTXUow0HobGAwLfF8eB
EizJqT0oIWhMLkaqJsXVMmOHCAE4E+DZimAjsn2eixvR8YDttY/J6kUdTsUt+pqp
QIZze++L5j4c+13fY7JR40XS3O3N1NtzhlII/F7USD+bSv5ics7CTMBWhUC8b5CH
TBDfP89Hze1FJQyTHK1Qk8Dy/o7OOm0yQ6YHwWg1l5UR0vAZm8nS3zHUuio/RxvW
GY0J3NRqjq0aYfaq7zyhVRTPeWfltZbMXm86EGCLDjAnMzPs3gsJXi0Qv7AncoIt
q4/CIQDlHbxD/5CvDFdFgmiu/LPWWTWmOdlxku6AdmfCRmFsB6Qi1r4so89Cum2J
FMOVXwQmCUHPGxuOWYnV2iI0VFa71qlBjfNzh9jVfYBrJxOgUgmAa9F5bZEGWTBM
vNP1KNGnHdguFYTWsfh17w6WaIV9sDLIsAG/Mn/rBKnKfCmHUbNVXrXr8YJODx9m
YbvBi24O4m4NIQWqN1vAlawJh0n3lBJxic1GG1E3kDPiMXDc8O/am7LtKzs5jx2U
tu4JZtpJ/mMii2W5A620TTbzZGRj5EmICRrSiJxica1Hw4iwQ867nFPUo+kAuJU2
iDxxJ+yXZ8yNpNWIoSvhbPk8Mj67icXx9lgnm/cM2yw3iAMtGCHa4JZb1gwAoTez
zlICLcrdPsrod65DTDRzxJUvcn5qTmDdjCqfu/U7WcsNAhlpq/UPYBcIFc9QoiO3
LD1O+ygbhJxSLtpuxACfg6wMePCXrbgdIdXbyIS+xh2nSPwMsSS3Dgbp4lu5X3mn
IFuhCTZbQmQ6JZv60r5Zv6OO5lkP8IGpFlVePF4QLDfaUMdSxLjx6Q5Up/IuIDjd
fOAsmnkR7qNHWbcqNevGP/pockcf2CAUKyxLMUdXfL7e2vvV4buUuVPhH8Wo4jY4
RuaHgrPe46JS+MqD6wGLgOTLtXQ2mjNIwGsj+IzqEsTpavDYZ47brADWwn7k88I3
mrMDunTE3o2hPMcYKAGvcxIcD7FMwSPkBdY37sQQ7yZrJhCe7QHm+WIKQXz+1C1x
FnZJFtvhmk0DTxD5F8KU1h8xaa8+ZTd20lnELqLDbwqb8T1Xcv2q9QIiMXRVoeMQ
gUt+z2A6EYT1gg6fXd17Z6t5gAF7Qt4SvFoBPhcw3BMFfNuZK+k6gn+Cgl8GWMlk
ku6aXjIcVbbD6hkoe95oLlvc5CveUQf7vv8xCojYjUZpNNC7gR1SZIzNqJdjRkJy
XSgDzASO8lob/Y6saRf5Ko9Ci+dhpAKs6cLozGvgQVMMkXmCumE50Z7/8WXEv3hd
00Y4b/+cxVHqaON2Fmk6x6FrvCK9nMc9bI5+bxoppm5s5DpI8BWvbKfbbS2PNDPL
OZZivwWlFk/Kpdr+MTh855ryWMU5+ZKfGmQdihgcCdlhuzhkdiYrdump2K7fmwbk
2B/fGnQFpQZY4Fo9VsvuRCAwJY8RG49P1ubqGrSRk58J/vU6dVqhSLHp6dBe237l
uZcvMg65qwaYLF8prCBg8vihK1XHH4i7N6Z7iU7OI9Kx8PyBg/O6E5Jvs/XVTlt8
5O+4QDS8mwXy1q2RW3dPLWtZLRcq0OE/pldC2IipiGJ3pGHMDlK4AxDjjxxGqYTs
+BJB1+Ie89x9WyqvdNpXncrzUaGvtdU6ij6glBurOsNw7BcXpNK+8+xvaR+2hODc
iqcEea/lblNVFzudzVtkX830vrBNyvRI040tltXIsMHN3N4SsTV0eLln8KNS28yt
xh1lBbPtFcc7fIxrW01gv9NzXaz7DRrqed8u+Hey46XYxSvgppsggSkhtNhdZPDg
GFFE5NlPevBDWRSsS54fuX16kGaOrRs5F+p1AY0T0GQi/LDhFrJ7xcwVNimigoDH
mmkyJoAzIBQoMIvJD1/CPkdDW9YUABm7x6bSN+8yFLapMXY8Oiu6cYOGAOxNsUff
24qccXDWM+mF99tGu0ryalR0igrzE+kU6ZEoY/w73C/9qGKuamwd9lFQXDyJcAL6
Nt1+1IWEi4V0aZ4vjrBNn9QlnQaIi0MjxRF2GZ91zeLXAicp6dvRNQWQ+fumT9pI
r7Xbz6ftO8blkgnNgJvO9kAwVd0fbvK9Mn35d/xq0zctOZr9niJDUdVRIP3x73Pf
F2zYiL6Zyqh22nVce5JaRgzWMS1yh78l/3k74L6vcV5WfS06knQru6onqtAu34N7
FqJlLKVSOJiDRo7Bw+qS5DG+PBdC44eO4u9KpUZakrz697t0GjtLL77Z7tXL/VdI
NI/w9eNHhoq7HmXddIdzkZNoRSxs2RxI63tMzALIP0gZkELk/dTKDqiyCRwPU0v0
sxNZUpG2nybF25EqGsRAdsOhix8dZe8VW04NGLoYMMI0Rx1bLBjCAtOM0ukfmXgW
b22eY3VFpFa8UHRvqQ2CWcsMaDMW5kJulz+bxNfY/9KrcaKoxU96ITwaLDiSBwXi
YDIFMEPxc6yDdj8c1kgdea7DHVvKJa6JncxBTH5dOWxdknHUZtml5JVTZfppreiZ
zOJQbRjibglSEG9biI+5/i1jO3p1nGcdMh7hus9ULDtDbaMh6FKjJS9La81PORyb
8/5dXflc8Ylbnbhxk6ajOQiRc7fIwvH7IWN3AbxPPSDAYLdrzX7AOXqT2XreLrgf
STjDi2vpoem0DfxTWjbl9TnP59gmy5xZyWlshnHUjBHx+eKB4WpHD+zza7JSokdt
3UC57fo2RGHEf7NScnZkDHMS+2e7azyUJsJvxanbLvNLS7viYsyayOAtNrLznXUi
F2+kWwtU7DuaNyJSoMlDsiS2IjswSYNi5Ca5nz4kjaf6Xtek0ii2TvDN4nkb605S
buGcz5yA8zvvd42OQO2WVIQ6D3rl+zJRmODtxDkIHdpqAt5vYh37wx+TkBAQr9YE
rR27CiJ9+G/xm+5tV41KyL+kSZpRuGYwb57vKNsGEThbACZjlpABlBldNbJbpT0N
xbFQHc2yUeutcypyhySKPN1Cl3jK0aC/+WDjbWZHMy3xLZTstXPolTrg/kB6Bwss
CERFVN5/23YCuIjtBhgobNd3wtTRry/oEUL1HSxe3qj4rB7S8jLMG/LuqkJlePbc
5UMB60Bbk8nO0xUDIYGyLFRnnOypEoZsEaz03Jes4ofFE7pSaj4zCeQZJa8ZHje7
vz0luN3d0mm9aN24WBMD97VJunJZFJL1/gaAPA6GjdFCgn3kkx4qzCrLo2jz9OzY
TMUBVPbdvJVDLbEWA/2iQ3BOQ2j5FpK8283caxBFi3R1Wa0qkvpsBqRzRbDdMNic
G30AcxohhVIN3Aik1bDhr4iyz4r2x5+1xrTTY7dbJUTmLJjmiVcpXDsufOIAe+fU
DW9TRi1PFjkt9IKSGWx74RNzB5PIH3a1k+GXaJh2o1Mha+re+55kPOni+yw/OsM/
N3BYQs6RJUjDApZ2LZpJ47058mCSVExFF6Py8n6f8b4Y0aciyT2XT5UhTskAEKTI
q5E3Shr1e14466pxzlfDshfh5ToHoH59G7p0fstSkhDodwOayljjyAN5O3bF3lzR
PINmsofkpvH9rt+BmEXXMrTl2rZ1A95fdN14I6n66C7AgNAoiqCYWXOVnQ8hOo58
5xFRCY9G+NDPblaBEByJOm1GihAaimUbkd6AijGLD+2GLpiDpp2UD8epAw/yyPn4
uTwCn0QdwJ8x5BN1fXTYrHpQye9yQ87Ns3I3rq+WVi4TKYiHleGWaw4yFC1xUFnh
Ya9sdmk8DrfVGYtZS+piHW0SrU6Nrmh99Z6a+mP5FSy9N51175AJCVupmbkwT8sv
D/QbH/QcnaR5hz0y3PpU0/KN9JtZUWnHl20xNJFbeob6lL0EkM0qmEaUzv8yDCdv
90i7999Bfdoj/qtklZOPLW+CuPvXc46bKSTFvhmB4OtlTXP0Ik6kJwz1okbQn+C/
2wF57t0MSUgGhFYmHyqIBxk1kS60eBvf4AsBXDQv3Dy1sKV4nbPE9vK8+PZpM03W
G0LMxr4bTRnu2h51jbElk7YDulX1zH2wxHAS7xI9tiXbp4bL5B9+lvuWbkRx62CD
SoTyLCgLIKQcAqxdvs63RyOdvuCVM8zhspwSrhRpZPUBu2FduN+wzXrBRf5y5Qg/
VkqyOFzDO59rdynGNqYC5uMwp59mlhn64vaFP2HN587hoG6LHbha4mNM7IAYx9SM
PqkHFtjrj002V9HwvnS81re9muRNXuXnH37tlEFEDb+EKWgorIrQSImZSbryfLVJ
1vudvUlKq9bdwV9oO/9TRvkVzVe/+ysbipFGiHIMb8GmbowOVpbYrWAp/3A2ETZd
6iCfzMojmvpshSR2mWLr4mg69FBm8gH6nK+HYoI3Ay9gMAKfxKsFSpOyQH29XPM6
B2qK8o6G67QuRoYayGocYqifPGgspKDupthJznRL7SSVg5gom63LqcGcNVUA92as
edaBRZ1YksTVrIuP1CU8j5nhM8SoY6B36eLYPm9YeTTpUUIwCZJtvQZ6/KyAsT3f
bh3HS50bz0oFwi39wQsVsRvvA4rgPTL4vcXPkd13lpFCakYD0VMB2aR3NdgpzMHj
xhOS+aEzFiKcNdkRcTWnetU9WQPfDfPI1eJ7hHiQLxqj92DMAM4Lo/kqPDuUCmm8
caQ+0M046xuOFjFzcBBPchrXuAYJui6zS+PjCouH8bKGhDAVvmbfK/apvDbrG7dr
bFiwf/PfTuseaU81GQ0fmFeBHu+F3a6u8jHdPQjn5n/G0lKQORAKZOlG8ck9tgSx
19UPd/OQv0yHkXmVBbNYgp1NPmiVoeQU4ppb/A9spEQVsmXiKO5x/sn/3mvt5SoM
zH3PZPSIDu0sEObp0gzsYs5UyTK1AWY1tCqqkziwo0qCv1fx1GGYdoMv1iqyytyz
VoR7WtjxOUtDl2O66sqVvEkKkUwnoo1/qq3rhwz7Hm94evjcFPH42bxUDgU9NC5D
UkOWB1Z0Ctkr/8cwK0jzsLiFMFsiWCsWsyqF1l9cQSr7TO23QGkZP1AxGgw1o1l6
LmiCPZYlxUs/KD3B5ef2E3FhRy2cUmmlTlpZOw5ihgNvcBgP+JskO4eS6qDvBl5k
ekyyn+T4DjMPiQEzBsiFScpFZ3qa1rkN8y0fVum7byARcfnXK11va6lgEw81CJ3/
3eWLtK5FbPqXJKVCjuixwtBpWvIVk9/YNj+oOae4S0ixi36GmSu74hpH1A71/5dS
kFZc1JKRWIP+B5z+KGJyw490auMlwHmAyjhJl+2DW1xjUFauXYIPB4T4EhAdjl+U
OFj1oug3bOm0V4g8Svkv1QgHI2nuclezXIJA8YV/4c6vwvTwzQetuASEJSZbyyLZ
mNsPPd57qfmlXFQw3dRAuQCP8W2Iz5fGLkZ28GOM1KYlJN8auQILURKMi0PFtINK
9tMLO+cyHplEWC/jAhKLDuqJCs1ZsnpkWrRPXfmvD7XmN4SGV1nhRMeGEGFiBzTW
FFe62vGHHX7AzE5p1xHZTJQ9oD+iHqdiUELZIKvYsyeFDEugCRO4aUsRpCPnj4R9
xnugVXE4o7EaZkVo7LoPlrN8hkvoxoHTQ+4MKdrceeYWv8R1olfs7QVo09mNM4bL
EKqnOVedPaaz0XdvvPIODwrt2CXrOXW7pNo6EGhrskyyyOaM7CM4VcxMrLqN4eDe
0EZMqp6Mp1SB2VeXVYCBQG2Px1CukvuTLgCE1ZkzN4xdMVm1H8YXPf4D12IseVqG
0dADU5+YwDDK93tz6Sqq2m9q9BSdnsMpzoHHQJbqd7nbHT3lsIji3cAyJz1i3iaP
K/ZCSNI1kRSpBosXnMeO1Q4SLWM+rNYb00+S6DLsV3nOkVtYHly7Nm4cNt8ChtY0
Td4U9oGqUziOnKw4sT6eUXkb2lXM0leK+/+EyNpvhtVYH/9gi2QXCSjDu2FPn46N
tetQS77lwkY6fbPlRQG7XME6pieRbQhQLzUyRNRLWa2rCLFHC7k79a2LHsv13nuw
H5VfOjsSH/1j3EhKlpjIAakQID4udWbu1uJQ1BABmCoQvz7d69TUb9Fu9cbG3MJo
1UiFrlYoxm72G91M5iRXBQGkFNk+DeC+GY7rlTCz/XB6p0QHeCh1axOlNl7l/mw5
cqsB3f8EfhbsoSqCI/Lk4534WoJSz80HnUV9xZ5H6FTkoaqJf7gCCRsBhLYyvPcI
HqMdYTkY+jyKt4zt9QLShuodqzggFXshKhdpj7isRGGXJaYAC1gYb94Y/GnHjF2R
wQMX/b61+icYaYaoKy7b2P7RuvWoRLwzQn7PwUA3ymiv4hlCqgjeXSI0WACirW3f
dy3MqfMdSfwPjs6wyxCQDuy/gXwXWLE9p/AS1+KSd8ILwXsz4G8pJK5jPs6CTRZX
4Try4fuWrsKnwFZrRGuAsGJ2ROjIMEXXVDHciM83a4fjNvnA2xaKXoDRaY6l65g4
xlo2O1KfmM4QmnQ7kW+Sq/44UGBltLQLp5kKkIgrQIXLCriKMQajBp0aQxOajOGf
dMvGIf65hVwH+SMM6/2oBhrOpXvaIhhDwReuoN7dSmO9Boq+ZDztDI2VJv1kOJyj
7Qocs6Bgz5zWF3IUFHQ01MCDcdSonS0nacIjYgcrurn3185D0D2pkhqrsUwPI+zk
1QvPTzWcuzOkCHONX1MZda45myFWU/XsA8uM3oO+8HJFdwB23Ak8Eo+oAv2Gw+xk
x2tZ69fiJlgcfMOlNfcG2nAhGZ4sNa9rDOOble6Xx5Hyv/IvNDbLCo8oPaulZBNQ
VqFXOb6xFhyoOsXVt0qF0udKnO/eUznqvQJhiKFQPLGPP1sWCuLNogNZOhxL8B8w
WezUdD7Tnu2wbNlfovsYaO7y5AtzD3uSxXpSO5LyfbkmsyJOorWVwnxeuIWd6fVL
Ptx21Th6WZOMweynl9+UQ9695BRiDtsI8Y1XwScaJxi8+AsNPKeSRJFACR+KUwrn
9QUS3rTKn1J95AfAFC1hJTgHIl6M5ary56K+3XcgJc1crIEF5nKxCKTp5ATLPOIl
Zgh4RxkPohvFIxBmhK8Mwx3I9YLgaVnpNoGf87visTSvp6HocVA9b2W1Uc9/IZMi
Cd2lnd5RYPwwkGKArhdhpCsTCbe36JRShDRB63Fqz3ZqLzx5g37PX7mbrB/VBLMx
lULPQhUyQc+k+0/qJg34AQNZgAzRCvO2KBjG1guB0du/t//TO9Y5kXfoyJc5i9l1
7IvHdv3trsSAXJWc+eaYqnRn0k6YKwbsJm7IZukG7Rg6QryNdKAw6YyHZlmZ3Ay9
6Ms7uQgDDMBpyTHg5DX7D/5QqqD1dyudFCgSoE/GNcAWEgEUSMnLKcCIjg/cyDEc
DgUyu/Dfd9e4mUkmeEAO2gpRm0hKRPFH0CUQCcwGLw7RlWlN6XyRPMAoFFKZjoHZ
x8uCSPuP/wDjYMl3FMnj3FB6U76rzPx0JI9UM9uNHGSTOn3YVj3+DHW6vSEO2hFw
UfnkeiF3q5ezt9KTS+Th9enYzWXSoIL9VpoiL6nmKvjbTYjXoEMi3QrX5fHz98i2
tZEU6EtrjJSgWb0xtH8MfL8dT299oB2Lzz9ynp1+IjWgn7VXWEvqBVp1lF6H4b8t
egqF+ZYwT1kLaSWnIJOrmpMIAkmQmmLxHOsiWM1lzUEyDSjrL/4zU2bWQ3IqyEQX
KOf9bvHcvThpmAOIYf93SyeujmjU3xrEHQx0RZwJxN4q/9/1ZTioOil2bO/PH2jK
OJU41t+Y7fHdZX6ovb41KkUpSbbUBrsrCxFLUWfS3+3G94mqGzojdGPVISGCt7V5
cKpw7vTqIwo3oaJGpVOLZrr7USEpsOo6YFzmrbfZXBINVWJcOoEtB1bJxrXUPDpi
xRrCpUR1oaWpXXicSl4S/d4mbuOU0mDvUR3DWZS6XuPMAUTXfaWUBvhSh6ysXPxI
laP9air6HJRjZcwEMABJAQCOO2jzMZgASfwf2iTPfGFv/NjSWHL03LlyiJ731WW8
klh7y/SsOQFSVrrUzHJxgZTbQmpBTWmE/B03mepWcI0k2aNb4RzFsLWtnK7NVeSK
2n7GbMQey1xFERJ3VA12QAdd9gO9xj2K30i/gvnmRr5/JbnCSvC904B1q8sYPUm0
Y8s3JfoYz1SI1PyV09e9Jr6p1ecAZ9MzYWVZuZgT1vGU0/TqQkibIJBBCd80yZrv
jumTHd5xGk5AZdb6HnJg6fgu0/tqCKbchAojK7N8m78PmCjPcrUIxMHC2PzIz9rH
XIx3EVUCr1wIYdHb+LvooL2k27dGLsBoZBXj4iy9A085dL11nULcm4jc/1KcT7Q5
KM+hM9UfffGwx3EO9r2kvqmDKDHPN8EfZBFZLXZZNZWIq2N0+eSk9c/0k2orja8D
BVD0mhciDxx8MODgMavM36oWiWnUTvVw9mviEdwcrLhWUKJcU0ijxt5TI1tFGR7U
W7mdyx/MlnzIUy3155g5OD00dY6jMNwoPyXzhcOJ5iCApVgLzVvjXk/VCe0VjE7K
UhMDRisWqEOfXjfn5JVVr3snrgFjfOuylPbCzlMGX+AbNheVHecI6oWxprkD+UmO
1A8L7LbUF0RpAqbEP2Atjj5gv5zG1wuji6lCqH6hGmxJCLg1NzhuU0djV/5Xv6Lb
vMRtg49Ig925+eOhjrSfvW0tUs7IYgHFPy2VUXeL8ZMVRQp3rVQyta1gu246Noq8
n7iAm7trTfcCn/YkMRDiwI+R3A8dJmCmDPA+kbcKkp8SRMgr4nZHFKKbIBtIkeJw
cIfBVgQKPaNTGhPEHGYiczum3chF8GbuHUEJ0PNHw06taBTRBkpOcXMMrrypiK2x
7+JVDW8v27LZ0SbSFJ88uSOSI+aeKEH7Sjys33zAcIkYK3+1GYEDmFKQYNBhwn1E
e27boA99hmiDOcNy2DDQQMpzJdpMs3YUq3hs0Ahd1CQgs7ZTte3lAAc6cTcvgCV7
MV5asmJ0IXCnGEPqO/pw3HDpqc32M2vfQd1xg8Rk6Ygo0SHB4g2nll2Us7g+BGiR
xhcY6krf9MdHnB3CUfWXBPuqADedmP+zDuGqJvuZcFIMp7rPm8Uk6uOjCXpaZXd1
3KXjp+fNtzL8LUOHzl88kbk+CqfvV5kovbJxaWdZxnwEmJtW1X0QiG/plyCdelL4
WdeKyVjUvOOeD55ie6aZTtpGyYz/j847zMLA/gnVzG2NJIWMb0qe5aY1cb/qnVIs
5Nw3Ha83jdjP9/Q+MuRFfrbUPEl6DiVLGt8oIFM/jMVTvmYS3BY36VNqdXijGAMW
kIAUSU8YMrRqPC7WmE4lfs1x4fnv2qCd7Eh82cC/rIyVDlJsEqsZJUFSUHYyPXeR
o+ZpdHa2MR8vbUHHXVCYmEQ+P+h2tXau/A+8+Kg003q8wBhMabg5f6cGaR5hyKGh
En9aRlYE59KYxvdXLWKDtU4rlg1FvKu9qqR8eM8fNAqI+zX3cpkRTCEWucM3/kwX
qivjwsO6N44umhuudwCqd3dvpqYC9JHUMaf8pz07JuhzMU4PwkZg2CME+rmmL53M
psThx8hF+K+TBg8SFvNyn/oHanYtPIEM4LR1wfVHGThcNnVejHxaCEotHsQBd4uP
W6R7zXfI1UsXeecTSiyMKUBnlb2BkC5mshdceMGij9zV2NTqQ/LlJ2K/VhO9vT8u
b8o/9WiE5jgDako/i5pCgQFqP4hPi8+OlxfYkav5IkfCOaET+q8sNVjGWewVjzdj
IO4slQL7BAYFNMevBsFcWDDzYB84D57r9LroYRmm2FPEeHiaKGGCYhorg2RYmH/D
kwkYYio2YzGFd2vlJ3OnISj67cJ8yh1uAWy+NFqNcnyKqDrvJG6wiQW9+gBB7q3M
lVpF9QUFbGZS4hCt+Xciy/FT+8D0Kb725NOWmAyvl0aAhrk8lHVzooLAWcViFGZs
zNnplRD0Lo6deI/6iZ7QttQxPHPE9h3G6TuPqMcj9JHvtx0h3Imeg/jMKOq4Y//p
sgtUWzUN+nP8L7rluz80a6ZlIb9wQVVCkdXpXqH24fbqK9jb1WLXb3bn2tt0jsLh
x8VVFYEHViG8JhrPUalx85dz8aeMfr+EbaCK8hVsTYQ2Spck/eIsMOaYHO5kdKde
9xz1B11U4ngNDIxChMFoxd8i1JJrh+v7Tghd4AmXPXzX3C01oEwgk6cMtH+pL8h1
Tf/4u7X7ixrrsoZDZWOLMPzaifWYCeO6x/eTKfPMfsFkNkDqqqh9YzjSrzm5/Bct
AEUYeTA+7pt0j99ySKjH9u+AxkUj0ktdr4o9PPkbVkIBQrK/V4E+tpT7yDB46NgR
pCTx8HWLY22ZR8HW5YNqXh9UElsPTJWBMHWQuQxsoxKVUVrruIgmLRLYfhA1GLNL
R8lhqNu4JbLktR5orktiHrHGORd9TwiIFNXclpJuCZOWslxJUOz4Bz+VURvQ/MI4
wdq+D/Xxxkq+cINPnJiitCZxqn1nSrfAAYGUPcgJBYRgJt4vG8lhE3sd9DfI214N
mgzGDrFAOyBlJqX+m4EYKuO/EvdSOcMs47bL2yxbVv2qFz5pt4e6eUXvrRhKPcgP
hCZ615weycz6aTLsaEX4jO5sXKsn0cOuDuFX5IuDfQnfPXRxWFdHu+hQqjw0Bfcu
xoub5MbRAI8zAUo6vUN+D5pIB4P428gc9vhxo1ZhQaNqDINZFyo0lrKeH7fNp2Ya
LknnJML6s6aBqRYS9jRBuQIKqYcGSn3BwRefua8cBI3YVf1bZkzHH2vm8OJkWPfA
5Rucyk8DPUjZmK0Zim5Hvpi5LNDrcJaqUBifr+cC+Ik7upSkSVu8ryZLVajHkpaX
lBUTlrTmk43naGJ0pNHt1pDVBwfBBUFsAkod+abMsI+QkyAiYcUGL3E8rq4Tjf/x
kyNpuYEKkGSojEVMuD/u0QREwPRI70Qe+C9qAXqYz0wnWlNptJ6qlRqsuxaj1qmv
mYTMkQaBYLwGk9WjSAA2h4So9qHAkkg7hCXD5NaMMQlP9yEuVQzld9lDQw8T83Yf
xOYfc4Qinch1Uy9rn7Ukqq+dD0eEX+BK1bOdaZgoaPXtm6BrKCH6Fl2FEJ20DPWo
J33MtJBp3+ndDSrnebl5K1atQZhRBz1sxr+pqk/a/0Hmd6rdpcg+NKsuLh9oRstV
/99XCH8pvb6Ye3yjLFd5jHg3KTaggKILX2Mca2Uo+RcjqSJSfFtGmV48+1xV66pa
E8NpY5JTtkL92gTfJ+DO3AXVftfseE9YRQPiNSrru8dV48+XAxLa4CJQs/YcX/N4
vaP5QO6Agwv+tVUskkce0inB/Xj9T2/gTRYkzboUV0+h3TEXgEHVJs9Ic/qCx4oX
K2RG/0AvFbZyQhMtYtF3l9ylY3DL30VSWoB37pDnfYYdp9zwn37ZhX7xKdxdNqWt
kC9fpch8U9nKnn2mrjehqtA6p33KSMA8iU672IO4kp1gOak15zsOuz2lxQ38mwwc
Mhh4UojJ3leKoeetHgkmiVlO+4aeG/zN/9/J3EuE2WOYs3pBG3hw6x/6GO8v27Tv
uVwF1Dmkfy8cpDIQbIrcVoM7R/wQg186KD8MbAHKOmVbleKBTfiYOY5q5GEheyuB
tnUyjSZ0vWUc9k4T1xvCULAIGiz2NmnUOYGPgPSs5Wqu4pqbCx9wJ7M+V8DoHsQ1
ZolQVU4Eue21tDAHqILDPKJ5BqAy0PxNRzB+qi3d2TyJ+stpZ3qAYo/3nfItB0bw
G13JgOY4W7aFF4KZelSKcbGEuc8FFfbHUugHhl3NCFc7uqbeqZEO+ZkoAy4ORWp6
fnbKX9+MF5RlLAW5ZwSZNoVDeuE6ydG+5ZNr+xx4pfrIZlZPUolipkbgdpdg9NpL
oLarXMfF3s6cR+mCyeBzkAH0xLaitqeVedXKqrdPgAEkCLbBYX2EgrRZA1eEoi2V
5FfV1O+We7IFRyvRaDVRH4zqio/vrhOgNJMXi59PL154r4r3JhiN71dymnehaYrp
2TPBg97ZN/rsmB4MYtULMn9hpckgYXQPqZCeMJYqVy8+1HN6szvsEywsRqrHB77g
3VnyGz3b6N/YcFjHlsB2rsoZm+idcSSIMnJW9bGxsLOlYLJtFHaXaGWoHOIb+PYx
EouxU6O4nqsGQ/HotIxCqlBJkU5WCApd+AH3NKHjZkb3HHagxADr9cOepoF00n2v
PVxtzz4a5C+2/bcBVjaPHXlAlMpGraZlN/v7od3poyqKTYyVsCi+oq1isobXKe6S
nJupDEOZa3zslOTEJkZf7f3Y+AcW6FXbn5p0RN3GZ1gg+icTKg2ZAIkxi0/aEDe4
JxX3BVVmnxFFU8voZe45GsKrh482akfNUDJsY5GJpO/8dEMCnx9AcxHPjmI58rvh
6J9Cl5RtUY41yworwsIe9/EheBKh9ItZ+Ee/0u6NC/BFQqWNXFUrLLw8EISDnZFA
SBSqrLez7QpQpda0yuDZh5KWh3dTY8H/lvUoKqV/upIMxUKOYJJTLtPDgaT+Mxwe
FswIVAu9IJbTmRlV9obsLpulM5BIBx8e9sJhYMLCJ/bEYryWB4NsQlmDfWys/W4O
OfD0hyRI6JH6Sy16Nro5ry1OYqi5fSh9XBXdpbZSrkQFt4vPluRdwitQeC5/ZO6o
kUgaQTe32xQiV/8ZXHXd/+1r1uR2ESZdHs1bWdXN5Y9qqPylGSYlG0Z5K+wcIboF
LsJit1R0B66Ch4pMYjt++8IMmtOGVVNRG7bUjpzPpbAb8V/+HrSBCPTDvl6MAebi
9XEx0M5uKH3gdlE9o7uQNkDU3zLXIwlhbAqT4+8A5nlL6czPjC4AsaSJekJ2H5HN
U7/VbZs3vpgaZygA66laDZB4M6QZBiln/T1NaTFHLRz0Xrf8DC60QGkjkPZeVLI/
7epJQAJTygaq84VZIIfSD7ZFpqi8Vvq1THjIxv8bZN8HYl5ggen0nsx1LES4XOS1
//sF19D1NaQkGKPXvuVCp9VqvjBCDdSTzUw3GYBaDfOP46nAwqaI6CmT2bj2v1sy
Pz+yDLMEBg7PRq4r5w12MW3/MOH7DAxVN7o5TF402Vm+1t5F0RTsSQ4QTe3UPNeW
IrnCCW3LhtEKNxpY6bd/kWelLoE9QK/dWoM9mVJpF4E7liwevHXlxijCf2QxbVlE
jxQCVGTDOG3gHeVUP8Gimix1Nj8xu3LAPBWEkfUibtVdjIv0ysQVGaEizfx0hXr0
cjuM5ZiFE3M4xVbLpgN3ZSbCKWKWB7YmVbQUmi3LM0pNRnSZem3v521cAT5Jjutl
6V6o+dLNG2fSImf08gwldlTIMVJTUjAtWsTb0Hh458mL2HvlYU8tstK0Ies5YuFl
iWNo+5tUCyjGH0mwIqjGPGSerJJgBSOd7fcrkoanK28sbQWWYPh6fYyrAB3FPmoP
exThFVBdQW/NWdb/RL4GEcbRDrpPqrOg6C1kLoyXu83iFHog8PiCGHAnIYM2Dshf
0SJyxGPa6wgxR1T6WoqOoVd+W8dNjf6V8j54E/jd5aSO7ngzDNu3885OPG3lxZhk
XYhF5/TZGnLufETutXGjVah3cb2HoNu6cSQEEAcQGXwkKHNP8WAx/sNS6DFYbiKZ
PNbh9X7Na0UZQ8odTLg8VPd7RuUjxGjfbOHC7vzReNGeFM+c0LvOVmUfPcerBsbH
wWbBaM5V1caKxHf9XZpQj0hGkpM6F9uivoz/XCoPIxAO9/7pvewAtOf+yWfNFgRh
yi1bsFeyTXDm7L+aKICGKPvDivPUlMdgX6OEEF3G9K6Sykgrh4aCn58gs28wY5s4
nu9vZEqPgP8gAOvMAeNUDKi8u9KhV1fQayTF51v7OdcIc4S2MGFupTp+LfqptTY/
L1hmdvmh7QjF64IEWS5kDZtyqi/fXB/1YEouFn3aJkJi8EhjjYs2y1p4OSLlNPVo
RDBHbRO3IGD0ay4HRbM2nZmFfxhAhM3mK7f55mgWAZDC6nqIY70Tk51PL0UcmHJv
6TUAwZc7RGMkg6VBNVgQkQv6yJFjJFle3Da3JfgVKa33fgU8XSTT9ZxLZpImQ/VI
PHM9556fjrr0XATaJnyvBiz79+5/6XCxQxo650+9XV9FBc0995agZA8kbmGP9H0L
m0uYGRdvycp7ZUzZmSATO5zdDxh/GV5FHsgjoXZVRDQVy/apFyXcdpSGyGI5gH7/
WG92R/0V9GaxW6BGHDk/dyvFrnlsieQXbeP0H1jV1NzKIvYw8YKjJc1jlmDCFzVq
hxSuoIxIPqcOfX2Y3g3oxRIE8eXtQYSk3MSMuqJTOlZBvbMRbx+CouBmS3GbVbfQ
0JUooiyyBGTR6ByTje7mqgRuiKKFIv9WLrPvoe5gZnoR4aWGtiTGsyfEkNjxpIAf
APHVDiJm/qaFjPS6ujLU1Y6z9111U8deH9LFKWF7rz4/1GgqenG000jF91RKjuaw
HMA61TQ6MkQao4by/a8V5nhu1chZr24ZdEkZJvKTByJqHEjE6vzK2/z2QIOGywKG
jOkylqZW0CjPNKnC0EuytGSAi9uT0EEBR+sfMih2lB81F0eSf0cM2qmN6WE/ZfG4
ws3xcP6U1OfW/r0ThMcJXgcoOAylZ5Kg9wKGzBWKQPS2aSahi99mX23UYIvm+UF1
rtv89AMt36eTRimSvXomnjNM6SwKG2mCpuoq1UpfzmZcOUE6DtTQt64tvDdr9cRg
/zquqP4mLc4eZ+buocGYXkKkBQV1TsU/QExDxJwCHmaihL91UjEUep3K9LhYkbH/
2P78pvvqFYhRhg3bLNscJWHhrKkZrxhcWhtfKpFLiMClkhpedAYEnlu0VSaWRHnb
oJLnpMbPMAN+id/5bvUTljOeB4wOSuqZJAxyoXM5ixa6+E43pqAs6QDxxyaRgbjM
N+rvyG363lkskdLbzlQAROpURbJk/8GdpviUfnVUMK16KxnyOuqojLlOQVdyUD4o
yy19f4eyNBdEK42nZoS9zhYXugbDel2Qss4vKteuL8vSp9kZs+Jh9PqJ/r5yg1nO
dE5mS0xP3zVk351suO7oILaMAoWYl+nTT7d6UpuDPCc52bIVOavlkU9UwMQLrazc
yuzNBSYOaZwEi/Rd+xhCmp8K5c72KhMIVv2d/XFAxM2kvZTXOXnId3QjaxGY6uXi
0wfaF5WchEDc0eQazQeTmgutyc1UvW6x9SYRPHtRlHi1br+6S85IH5yQ2y0Q1lZ1
yhnrudp2ZSno+Gnb3PVcpUOj3zJhrqZ57Qizw63rl7cMRO5eu0Lxbt0rsd6ksy+n
Jh/YUjTbcZ5VRdSwSgWMo5Qi9b7gcCtCUodCYb0Q4Y8SYK/2ekUssFZnbo5YkftY
2tfM9C4fYOHlTiBPvVXQjuedphelpGKI25RAhBnJIcyTLu4WUwK3GFs+TqhQytFD
49HfODLrZUJxr8ceISEWVieVJcw87jAlLXDBglFZhXXQyAo2BS8j9BgSaZQI28am
CG7P5KKrHHrim5MfQGyA5BchL0jdJ5fR72qlYP3hmKOn/iSnc/NAKDjI0oZamJld
MpukJK82Wa0BAb6ohny8KJ91978xa7c2hYZfwbCxfSxmcbv/VWT+2iDCYOsXLc9Z
d1w+OtQkdLB2oQrESxeUoGPe+0nTauCn9aT4gSThCfDEpHrEEnOcm+9SX0XF+/xb
IJ0yK/x1w5Yw1+vxs0QMpy0LirAcVU8i3D7yq+SXgBgKXOAyyJ6blImL13sd4dJW
aRj9CNBW+gZVOK5fSGvv5ekz0O83RDHWKS8dLWfnTRZnr1dsELlvsHrfL/hrQpCA
m85JLb6sELNBAoTzstJx333UYeJJPDxg+qLOqB5Wro9XyADarp+7gKJukv0idCok
g3iYqPToutm02xg313r3SIAEuXXsAD9yeky/CFLMlFyjFWNdAqMNFf1ppe4s9u3q
zHlp1xHud9cXzLUeCPCYzo5gtgCds73QlTwqxS9z92xStiUs8ViDvipkcPKQK064
zFXnqb0FG9aBDYetjRBuXM5UNFlF9C6Ti6+ck1Wdbf21oCuOk4JIoWukIsM2KrQV
XjFDMjzuIj+/pWa6fOmNFp7hRErChjSfwiYAHs0R/a9UGA+UpMdG2eHR1+Njhef/
M93KnOPGpkbE4udxq7AcJ01TlsJPD+XqhB3kqQqQ/n6F9hk+L/BabRYlpF0KKWil
uR2NeCJblBNBgWtIDRo1xBykt0e5rpbwKjdVSsYcGWhlz4eFGd4CyjCSLFmJCrOV
Zal1YpcihO6j7raXEaifAmRAl+tM0ra2iuWgZnceidWdT4dmne6p8IYAB/kTc2J3
dP7VfMDD2EzNNy+jAtpZdt1/z0I5cWqmIOH0dkk1UNgEyTi9Pv+Tnk/NyBEW8oVN
XhXypAAdCuhTXiXhXwA4VgEmSs3UdqaDpwNUskAUC4v+n3Mc9UT6EOQWQ8JL4y61
ZRlRWPOo+l67g0kqOyXn0h4a8PfvQ38ANP7YWeAKl8hFTOQoX0niNgEmB0hFP6f+
1pV47cEur7e9kA9dLef/uzEtRRS/6JPVTLEpcdMha9X2JbhmQzYOSEFlGWxCPTdO
mvhzb2auZ3FAEmC/VyuZqCwmVV/EHrXFnTEr3k71vtmDA5jT0HGVBvIYND00KTYN
dYnrWUIJ3yyjkokzHkwEt1R4YIDG/grGK7Bn/byhbVm2hM6OifDC4vJBIQrPVNAS
DIS9uP+XhMJMq402QtLpvGEG5z039r8FEAS/TrmfERX8KpowzqKQ341zEnnG0MHn
5CmnVacx5pALR94/j5GxfF9PUJ5zOoAIBVOkcMBkWaha6fAMKlpqlnQj1QkZu2Gt
WNJb0Eyb8LT18mR/c9MAeTFdKC4hHNgujQE62rog3oi5U+1Ifllb/w4VwfAPbTuG
UgrTkZ0QqvQaQk7rPGd3xAxP4/Q/qbhGXt2zQMa/Og0+US8AqUtricYtvFfCveTE
bFgpnIx6wbn+V2ofElLh1in9n9BUsmVs+pIl6JO3bW1i30eMrW9Mq7evc1nclD07
SQazWswoN3VnjMj8T+hd3gO04DcMfHuGA9m1kCf9496HTxV2Ae7yuoiwjisU6vj0
Qwrev7YNRgp0u8jku455OyuqvhZSlW+QAODi5GphNlV/VWbJvrriOq61JtUwK4GU
adGA6W5twmDBBBLr4PbZxYsR9DvJdSztHu0pJELbuCc1Kdq1nP8oCEZsJSW502XF
fSBKXQirBs6wxUwJasuvvH0SH7aW0d41DDm7qdfB1fPnFOUIpe7DfiHaGpMgJVnv
t8ncmnuKFTmcAHt+eRI5s5MWtHRsxnf+MglngbQbjZ8umLXAJv4aIG1wlo4IOvtN
DR6/A0hHSINxNxh5zIuq8u++n0e/gDNisJC5dkuVsachqWsXZccOytA3h1FfyZMb
sHnCiMIMHHt9lW1S8MhEULIRiqBpAWVDkJf1YYIuC25DHBTHtz0rM9VqCehAXym3
ycQxJdaSmzE7pBnAfnl+2zc3WdSZVS54oke3DDuyXdrHhwnvHi7OoNFJ0BOq/4MX
yG5XNgXl1LqyDml9Z9OWGWVFF53W3vOLboV0TesOToHH/MXJ8ze5ntDLpJAV//Gu
QH4tvCNKVG/mvd21kWNTe8IkxAgrM6OLqH9smM5oBT7Nt63VyBuRRYxvP3sKn9IA
dMNdnXXjI5hpL1QLV4qiS5QGxFMPgRWkzxUA6ReMxFxCgZYQEe4/dNH+Fd/l2ImC
W5W3FR/MFfuje8yLEwiwzB6utedjg1pJTssLwIck90HOApkqhTh67K8P3JA0YyWE
bdTtv/ufHlF1dSaWWh9G3rf7oWRieBXxfEdhMLfrVRZaeKYVelaXQineIg2vqqCe
37Tgux/P3ANS+6TuRyfpK98DkpTVs6bTauTl0C2ng0YWWMtayaAKWspWBMgskirU
ipy6yhwsEQrT6l8RHkpiXLi98R3PMFY3MZr8Iyukka9OmlYVM7bWKSTO2KnrwXv0
pm0Hy9d5PFHqO1r5hq/COl/Ib394CYdFSs7GDKIPjTzCK+E9aYOvw8z9xVRMvOuH
FunJtqi1K/pGYeth09i8RfnvYqWMNv5gOMAukZoykS/E9I3IR2EdEmzI959q/Yr0
3SovaR8saQnmfodM7tusEdehngBU+OQaNWPSJwn7SdrjqfqEPfLd/Qspp3IFuonP
I1/gq4gdYvDBrjxxYFhr3mFjnuIHgKvANgg9f1gdepd7HGkGuUvdvvQAThh5YEIz
3+svQcEWpLAu6A8YM3abMzNJdheC2XrYsvihqxyFHBrBP6UdrIjTg0aAx+nAEd0s
eS4Ak7bQq5nWrGUL4RORqw8h2r+629u6QJpDM1bbi4FN8PhSqHWGCFrlQFFsWOG6
onrDTPc5hOeIfB0EWxPoPYdO1Le8AZPQludoQimtYy/+6Jfypo5eiXLBMmwxrNPu
1LGAbGfn5S3ksNMJE5CRuMiNQbGcgcJs7apieOaTR9P5NFko3bBQ7y1is9Drkj+O
QhW6zft76o11iNRSWJGvYUlKu22EBa+AwZL/b9LoR+KIKMJUln5QxSsCiabMleCX
joZOlv2y2QPFjb18vkVCqfIP0N4hpUv/QqX68sT8lBe6Z3RnOJgucwrgVaF3sQpy
LttHan4oX8zxPM+sLhIQyxkUxTtbGyltQaeFDp3JabzYd5SA29JhAGxI489JVO8r
TDjpoMWV10ab/q2yxLiWMotxt6zM44MARD464nxk95KBfWR5M2cHAe5QgR773e4F
c7761/npvbP2XrPYwVy7nMFYD5FEYxB17fzLK9TKxfJMcjuTPaQDmM/JQH2y+r2u
gKq7Am6CmVTECSIbJ/5klOyq9hqzHkn3vWIOvVKlHmt7w1u4EBtC94Kx8cdcpM8c
H7rMARpQWcR5WFjQnrLWX/4xpet9hsMOXII8cjUt+4TzJ83LYU7d6LFvw7Vw3DhN
G5dP3gjEVdcYpYp9ymhSz7Gd3cRNbvn7Rciaqt7tcGSxhdEmStq//VhEAtxMT5Qo
ySOw6YfIdOgv6A5Pf+pLQ7UNFq7xnyT8moiogJTWJrtVy1nSjMvvuEdhpmjcfXKK
jRoSTGnHPopACmoZv774HllTDH9y8FcWBrBOwakHsINbMBg6SiTbMzdKbEnr73JG
4HstjLJf9nRhN/1Mz5Bb6gGqgc2d5Q8mPz1dLQTAQ7P+10BnM460XQ2oP11AWm4E
F9BE8vG0VjLYczMePZenwkUYq4kt3hQGhDE0GZQjQxhkl4DEKAMt2RqDxSMkQ9lX
E+aMCaXz7sC/k2w2Z965H/QXrGzBIoBPJVQHojTuAxv59AVYkVbKHZ3TLtr0f8H7
XHbm1cpzpjWcx0OIIEqji3IwcgN9HiaY8Z5yoHROwb84jY7GFiBNrC2oqXFpJiV3
Ig01xIGGdIn8Ioqaf7yXUji5EEXcxx5K4EVbfaBaFKlw/P/10sXyXwOy8TO9XJ5I
PRE8pMe1qtQ1ujSAx2aOs0qIw0QsQN4Nu4LGGPnoyVKM/H5F1e/eN9xdQpixZRmC
e+5gbC8a3TLGZ5tNyak2YV5B7hC+AgZtJHyTLUP+K7Dayvm7SoPqN7GT3LniDpF3
qykmk7Lvxv3rZSxgPbk4gBNrLwHnulxNriu2h5hdEdXFVnGYx7v/Ro4q6fUItpfY
Peq7lotm/aJvy2TFwePw07BC1sFHz2hLeRjqq/wG2sELpLF8afjNAjTDYBvR7Daf
Qh2R0Ow92RDrMxncaOXfu/yXcQPjgnrzsgxuSsPmbwqszpumcCyKTyOOqCahLANQ
8bfFHG5zTOYErfNacHnKJwiX8vTbkT9DZ4nnje3eSCcuL5vCysceOIUGrUGYCSdu
MnfeRljAKYQLlqjXxyK682s+LjPMCZrEKf+MM+55aZFOLLgQRXqSO2R39ZmgpE22
ocd3xeEPfDr215OCWJu2YGpHwJBYrLRzdhaHjg2A13/83G95IqDguNQJ+9wrJ/3y
TOj2ypG26HIm5Zx+NavsJ6wdlYh1K25pX7Ra8H7AlIEq9XilpJWZ9RaMIJrAkfau
TlTQv+IbZxlHUwiSuL6o25ASO6GUOMfU222NCEpCA7X87ga8osWhet/FPvXtUEOl
hIhL/vQDTh1sHxZzzJV2LUP4bB2qjKXpeHofZxec2ypQ0WT9coHMbcWMez42MIdY
2VLntbUA/5xZvuORZlKg4z7Z9HYsOLf7yNoXWEzMkHsYr9xn+TabP7Mvh9qPgf9j
LxRQZkqwWtphCjs0aAwYGIENdCye16emTj9pH6/SqO222JDRVN8k/+9OMqtzgeyO
d05PP1I9YR+d/uezKs+Y5fhLN/QNZBgF7dIrpN8tCm+N+IjB5wCaq3NkNL+FgyW5
dm1rVaJMtmhA7qfgqmjFo+sng2DMcRu1cZqSv6ffsdR+3CUS063B77O7JQvU+VEr
FDWur0ReqjzCQwKp8V9xx49EPXkk1P0MBN6Q1Wf5sS7fv0zcgS5CnwepPrY2Z6R4
jgyDtT+9NmveGmrvNFn3amIbwml67ZYmVORFjqWsDoIAb+VzEItjKPGvE7b4oNQ4
2Stt5tvAP5CvTDGoOqbyI9pgHHYGJVOMiFyzq5Pz4897TnqOTyMuMftzKta0uG7S
1VCqN82QZQpGWsDJ9kIDFV1Z/xV4aqNJvq7NQlrO+hiN6/t7UJ6U4I+azw/1njUh
rcUJjKU6Pa0YsgFcp9xljPUsN/J10mrsh7UNFZ+phmFSMffgj3rNDU2P09P98LCK
W4SNIoTCNXbyppmqPRCrX6SeR/7nuPrQ4zggdh4WCJOQmXRDp/lODHUYiGxuB3Si
IsZ8OQauXSkz5iGsxM8ObOJn/qQpIuq6LFGKj5PdyQmxMkQKuxdKqxFQ3i+T/8Js
wgZYcU6gTp/PDHMzzjIXdVG6r1G4auaC86Q2n5HgXggBRIPQt45y/kKKNiqFZ4Fl
PuBJZbfNsj6zI50Ce7WhHMJmGRe5+DqRV2Y+qZV6pdGw2xiH5g5epc1sPm1tBZfo
Znwgq06FfNzRFzwiKgz+9K4M+r+2o5OQ1WIscLNU7qa9VcW4w34JkIxY9eXSlXjT
MiUzNj2vvm9rTuh3suIN/uvagiELpiLYzJ3ofV15wUqqaXDwbwTPgNCkf07m9+K2
C4iWzZfV1MfIY+WX14w6qbyEKCw0N4bzxe2mXUqzxe0EauOSlU/xF1u+uNxT+rhz
D0LNurWjxwh0c430agXA2p+kP5znqtTG3yweL61FSoLkclMng/DiEBHEuHljBjxG
eE/UDvzKJ/vSjNirGFA5NxQkZTRTexSrVAr3vB2zDG/bPX3L7Sl1pi9Na8zEJ23/
YxU6EGHaAExrQrXTSoNVBAU55xEOa6VvqiahyvOrPNiVDiGGEdGKZTYFj4dmOhw3
PtqSCbH5mJJCIApD+IJ6WIUdS3FBUgx9Hs55v83EBFYk9dNCJpfPtpm/mquy7gJW
PZCiBGDlg6OXMmh+4PjCpPKiwFrHN7iiiaJJRXWk4PDZKSdNOYH+Dt/rxTFBETUz
1BS836YIw32s2bLvyIZOIKYwY/CwtxMc6kShkTbi95FNBWXeSo8He7rl4XoXLWLo
hU2NIkW746L8Lk/DVyLZoI5aaUkmBXaU/xhflRn7Vh3E9aRF2LhGxRLN4umzO6S1
DRAtzN/vUM33LvUMgKCwGo6iOAQLo8Od77+4VAMpEAYx1ogXRns7L8jhFYRHXrne
M9F5YJde4t7uRxL04D80bBO6u6VtQwY2BWXALrB9FLggW1RLsfKIhEJ+X8S1QawR
iCShCA72vRzG+LTlBJYiUCzLxqu+vTWfhs5amICVmcfS7dmZTr3SxNHnvWGW+U+J
UUFnCWH1tUy1J7rOhuVK19fHMw3lign11z2Q7TNo/g2Co//6pXv/sq+9GGmpoZV1
ME/wwp6hVXRoQMaIaQCOOR7PeSmVqEok253Ug3kGCQvREEO4sqFsud0I3YxlLkxn
gfuKUK3Ev6NBtmm5Q7D8kzYhaItkf2A40/Z7As85LgzZRpEPzCENGNl+stVEJaZ+
hi3lzyfNi22CZZUIdzTZdJEgnIRPpeQZ0mLesyFeGskQY6x7UBjt9uj7gJ6JY3HY
BUaTymg1u/4XfQAjghcEvtoqD116P/YMNKbnhPwCwa/9nPecNVGJNOmrynJp2eHN
me+Fn8t1GreksccVJZkO2BKkl5v0USW/loR1byh4P/nCIZ7n/7DFM3/9GK7VPIGl
uoo7t8plrOP9Atl4ZwyUZjLq3TfL+d2uf/qlqMJa2PrKLKOp6Rp6mHDTh7nSVDO2
eyKzrl0FaG3UnM62QF3k6i53cFkuO0A2/6UxOTRRK9nL5ULIcfncF4+t7V6z54zw
cQlIDvZ/O5nooTOKR21wJbfiLE8Mgp1Nv9puARwRVqp3hPSeGUlFXZ3zQD4mU9Ab
KPOADq7OodZnNXnNK95kDiElVizV2HBKm6qKpqJIzKxszwHdAk+wCYA1UGKftkjY
0SaZzKeGsLqQlxzUXNI03FnWSt86rCFwuKjLTbYIP1oBRZ2DQw3PJCyqFr5am0ta
Hl3WER9HGRdVz1kC025GBH+RNwdTN/Kh4uVzajmTpVibIFZT5v0dWk1APKcVj6Ev
nTdpbLNQ3iQEZoHm57FHXjGwhhjwe3NBacu1lHGh0aslhvkD6uLlsA5tT3aRx6bP
+d76p6legwiWUofbtwfbUPtXbWHHKH5ciqd0p9cWBP0lVlSJf24I39mUEdoSVqqs
efKvnXvIyEe29GjhSCBqZcbR3sjgHkGAnaNoB4ARL00gXhfll/KVpkzj/f5SMxh4
u3QHYDLhSjKSXgS1/DOD0Nqot1j2abUQMeHLhPkhapUPoXB1UdQGAAs5TExURjMx
Mxq+wonZpeJ4PqRdx6/YJRq1ufwfsHmBXtIDWlaWBSqtV/jza20ZMxH1q9YghJk9
lkHzou5SVz8CCjXPpKfRHyPCaL2p8Fw7N1/aILTrNe7bXebeuPYsrhfB8ONLgPSn
/l8r/1uj6KP1eO9WzxgL8EhHhK3vQxZ7rVgNzc9FSOmqJ+VSBndTyH4YN9MZI35g
XMKOoT2Q5Ay+kUwv7rCwLT+E+XqyYyTxMMvCC7ExBvtEu+HBGYSX1iT8+FmETiFR
vXSkL4PYh09UkrpcIbsDHSUoi4imoaZMRHD+rhLDan4wr/FYNg8ED3J7AzuI5bMO
e/czPkE/+tctK3rs2Vsnp2hyntAruUjWtP8+xAy8rJ/yVrfw1i9xnlDwXMxrEhwl
UYng7ZKrznI71I5B6CbWAvjF9X9xB3Z15cz/ZSmcVc+83TVKjdhIk6iaQjgN4jJA
yav5flSBu6S3RIG+95wfl5+onoT8Ck7szmm5mW2jaBGbRn2yjcN2ul6haWkga0SU
bLuQ6GpZNQQa5x3Z08zOPt9YFl8TRXlzonnRXwUlby5AdxfzfNjmQBoFCq2ykcSd
4CThTkworMc2so4D0GNGluSKBUPiATRi/gpKtoKKslrM0mRpIhiiR2p4GitcBzFX
dQHC4eyTsVVgleJv8qKshoX4+ugRMP7O5kU5Q/1x5mv4dqRWTCxELBUhLGVtGbwM
SluQYEBzl3B5mH8+dbcajz+xRQa1dFcY/6P/Ini3Pt+ljV2QPi9ea2oxLs4XetNp
oQOCHhEFWuLAMDwdvwJAVoVlBBc2VU1xNeb/XluoodbgPv3++IU+YpiG2te8JIB9
XFjDWIzIs99jVw6JUkWvGnaH+e5/7otE0pGUlhh/Qt4wnupaHBuRFY8Ta1NYlnSH
5ZbtvGdPev2do/GYLEuxP7XLgNa44kajXwhoDCXlwVPq2Oae6lhxKDZCyhm2byuL
tvjeom8SrKakvdDDSyTwJvoaeZcaAyHYZApxbZ3QzMwkAgw7xxM4HuYnfqJc2O3q
gFuHLoyT/btLfXrFx969WbeVY3T5iok5cyVj7fDV1KXSb08wabxLreCoO+/0x1Ax
XaXT/PWCcIvmaz8pS3mXSZXQq06MZk7l6G9769Nz0+011h3FxDZfab754GHmx8v2
t2zRa72QIHqUSf0I2K6m7wNesieOe6l/hZAicmHtLChjnjiK0cK02YSj5yy7lFel
J048PTo2/rZCl5LQHvHjCILykTocm67h9MfuX3MmIcFIr9xTZsAJI0uKWGnXVVmf
01I3GOX7DE4JVjjILJPC1XMgnRKX/uL1zG9/29DYuQTxXM50wKrQZD9nXs3fHf2a
p8dzWVoRHVmBrzHvPR0pxMEzVCqaO3o4ohONGObkzQlawl7X0+D+9F/mkc+XZVPI
Ix+5yCH28e/RGQGUzUL67hrcAG+uXih5P4ciqGzGtMFu3Kgw1BxtHIkQHOmSS0XJ
4R2hOST1tcVCZWpkTXcC6yCkOY4Vhuy6d4keKLCGDAM1bK3jRUl0IP9kntgaPWbl
O4XpMTqyoDJ5k+oTs9XEdYmXgE+XI2J3Jo5zVU2UtU4mvjn/OOjot+GsqjCY4g4k
5wDhBD2Ot5LXToTqOk1Lz+rXFlunTIaeikqn6+gGkmT1rd7kXpxZKgZeUXRzupC5
He3ZvZIlysj/QPLbn8T1bhPrKnDlyNfsxI8cwJ12h0Wq81d+LdTelCCYq1qpiHi+
eUbHPPVGMBRIWsy5F9xs5bQoqpooSLjYuZtXH2CjgOyRs2snHM8UsuPo7LNdEveN
CGiKKcqIG/wyrSLpr43fklyzQ8GxQNdE6D9PqCk6aBByXFc7zrQKr4wUNHJOkNCO
dK/at6sTwflRCUDTVH9kRAdUi4FX8bSu+kM/kos/wcJqjr6XhTwyZcgitC5NKbJ6
hR3un1mykv7C9S/RRo8wQRfwND3auaJv12eaTKUiqH5dX917gBN7Gv6fnZAEekJc
RtGcpGeksj0Ktdowt7hphE8MyFOGXaPRveq7uVbkMyQwws7dUmhysnSOP55rFG85
P92H+C4LhwMQdHtlebIhrln7KlIhEZMxJhTZpWVkIDHZSFEMUv/PWOL4Q14XaPYk
Svvu6DzedfHheSDAxsPZw8kyhuz0LgaCJmLaXG8I8IMpOboGs8Bu6GgqRJQa9i87
r8//RijwDszngs5pvbySqxlBl+qTNh0h9UfotGFxu5hKSGCVasw1kGQi2s1RmiUs
4YtpHw5olGnu1oclZtdyRrGiFExNmY8mhce+enZ5q1HYula+KbGUARUv0S5boB82
LW9nSNYXBsca7ZnxXo9Tx+14/X9wS9kvlTm/o8gIzTKwfRz0jTApOCTAB14WeGMr
tzo1eUy0YnEoUVNDWSUwkuOLh4F6wLiOB3STchNXEYtug/aVqrOPoKpk6NLq+e8r
gWlKWXesdGDt96l2mrCpDcdTVhxhj7nK33HmMi7DyWeWN/M8Z0Cg1yo/VKQeZXEJ
YNVAM65Y7OkIbCD1UlH5klSf++RmSzUQuUi8Q4B1r8xonyTZKPQ9sYLiPV5BrXFU
iX6K+3uYgLbzvkvnsoSferLW0ekqEUnRE0o712SLwEl4S3L9OVsn4GiJKhmlLKRs
uWhZCbht1ZEwJeDl2QfPtBrCE6EOjacinUumg+DT09I9ZghrXwKvTuW1SEzypEPB
H+pOFE1mawfN/W/1OLcVQmA0ntT/NfKEwf2fMzFJxnO1gIlZbA+YzhzyQ0pnHpYX
4iKxnr/rfXqR39fplUZmBIGgdBB+fGDDoZ1YcqH2sng1quLThJfm4/XClzMbKPWE
MSVVIwoKg1SZ0T5MYb+Rjea1p9CoziWAbO9f36shMxyNsHx5ICk4A+ctn2stgWsu
lGFEGjEF2kuyQVKi4ZYBXOmMc6A4E3rwhXyUVIX25W6joIO1R4A3GpXU08rfZ+sE
R8j45FfPrPovLsRxMz1fCWRn7ebYiSN/0U0ddLaI2j3SJL5BqQRRjk0ZstEYhCVl
KTwxzDnwaXEDKysvogalN2EUmsx/pFfR7vxizViKi4SORDUkDTwgEOVWPoYTT1s+
I2cbLzmEKE8GVcRBkW6yGLt8UjYDIDHOOqXQXGcOuuf3Mx2AxlJoPSlacKIdI0fg
FJxsEo/Kl0cvtAG0uwSoJJeb1qJmJCyL767ndLD+JLNPrMcVUn7V6x7Ac/TGUEWN
1hyRQ30uqkmsmZdLJiFkPkIqruIyuSWlb7SxFq+xxO0r6SqcFFWD9PJt4KQH+2zq
f2T7FMlGBVd6N6V0vEDJr72MX7NR+nM/R9/URc8WBypUKY1AMw70wWGZd+qcwz3m
63KCcUDNXIWJ3YdCVh5iA3a1icyFvz8cYX1o3BrkEFQCJV/0sZtCqqYHaGv2xPah
A7OVJHlpRn0eh+O0g74YBdX9rIqNYeMQNJRWckIR4cieXZtn2yjsXmupjPMiJiA5
eV4WCzstkD5goVrli69iv765nsyvw0PL1tdOPLEoIKm6xfpsZ/wD9bWIx3IGZT0Z
GME7SmGALe9WwlMqPg3CN2pdcg53eMNLqEPM9IJ8LEAjrkOoT61UkQsDneTBQhqS
2DSRrtzYvLVzdeq1YTut3zZdmCA/QiJjY64+6hmWc8AzyZ+uOgjirfHfqRcO2sGq
ZK8FCJ1zh2krEeXSxGKeeO4NBObWtTOneIRYs+YvuqoM4VCmvUczoeHyOkW5B1gH
ENw30e0G+1Fk2iDzGu4xed5ZrjUQohaUZ/QXRhUR19mKeSEnl0IVMT1s/7OJ8MQt
EigBcR7Lt+jNtBNOyXAlpC3KK4G4O9Avk01Ta4lKac2JvelxrkjHH0xeUYgQ05OR
kI81FsfGYw3r77IsxoncfftBWzhCtPF9mV4+o/TI7d5xwhmTIOFv1y/1gSVgEVrI
K5Kl9xvk8mzupDrTtHXXBctdF0LfStMUISk0hkIrn1oYNnsZlMY/uJj0mMQgqXO2
bv/bxX0lfd+n1XLGB99GiovKVTAOOTXrHTben0hDAffdgW2IGOaPCJWZwZFTg0/D
oiQ89x7qExqFRye4A2Gvbf1vWypVWSVXzCMAGuXIA2/mT1fujds69OSWkSvPkV88
BAFqGttRbPR24gy/PjDHrz2qKgU2cmJi33wHkoGnlT4qkE5mEcQoyL9txx4tPkVH
/tw8BuI8BdXKQMvb4HJPcE860UGf+9pyjg3lZNOT2vMiT8zwSOf0xCyB+2lw/wBR
TDOWY4QNdBUSg6YFIYOP/BmPCkAFgQf/SAt3AN8Fsd9f696Y3OEd3i/4nbNoxezp
QxZFKlTZ8IkXpX7pYcrD8X39/mVdIUYiP8fx7mn5gE82fnS5W86B5UX1WgH6UGg6
FN74lvK0qgvfUoFwOcDBaE+ETwdjmsKv8fh8VFvaP5uRR/ckIrmjRa2rRVn10XnZ
eMWk8Mo+txOKKUj51zrSdy8mNas51gHAtKrQLxUyGB8KOd8G9TvgqNnJvV29K1hX
Wj/4VHADOVQlqDGWsEm7LTpmzETh2BJHtYXOaqnOXIpfhT/pOS2wxHnymHYOfZDq
MSrxRThE4Av5ww/RjfD0EzG5U/qz3LZb/XFMGWxE65cinGTx55ldpQRuVoG0UHuD
7UyVBeJFDzwZUHrFmPpajBr16fn+GbXaUJ+FWAveO1WTEL3TT79/wgX9ZIts1jN9
yv2ggkryVnS90bAkYlJ1n+nkeklzwnN1rL694sHuhYXhzlSCk88htLW71Q15iZgZ
UW9wO+fp+d5z61FsRCLIIc456QW2ApJw3FiiiEfHEwPjQSjd/94yN5mYfQ6fEFe6
ccLZcmMPe+Qxq4rZii5Fdkoud/2a6XgfsRySDs4E5u63nIcObTzU7uLgKOnAt/DG
2H4hWHHgJtNKymmuexg/ThDKqjS4ph1t8ylJuTgrGS3eAgqM/2KwBeOe9rfD8qsP
FckgUKszaHLIiPyxpquzLB4hketjeIrm3LibrGt/Lm9h07hWQXh5rBkqvwy4vVrr
F4CI8ZfwPMwUm8MiZS+6+pbBw5MdyJxTP3Br4Xsc4JGSP1D3ph6jsNKaDJai5MJo
yQiEwHq2GxJMJgwK44dB4f4U59d6ob/jD3bVoUHGEOicZzFwNFeEKHzN4l6rdM0k
4d3c2on1Wj2YpHC/Tjzzp4A7gk0rq1+fX0EKons58043pM5z0h/27OnPSPAYHJS1
HyM7kezXrJzkJuScBKkqV6FzN4tReppSOQJPV7zU/UVQA2OLiIsoeULWjTTWTskO
nLluBezt67Uu1fvCkAwDfAHdUFt2dzM1qkwLFNcQDchxAR1zSF7Gknd9t4tDCBLY
HzMaelCTvQh4XF/ryxrNSSNe7lmLsHsm79Zplrusw/VR8HhEV4KyTdst9kzyrTEK
W2Q5inUokD/FvWJ/Arc0kfGONWbobLHeFRZl0VRHXngH9qEFJDjGByGjYfB7PWQw
ZoGkyTRlt1d0OGZLaYD0Bcj1+N1cdjbNnhTe5MYgMqkjb6OiHovbbc6VN44nuEhi
wyCqZN6lO+G7T0n5HKa6f147orKuzfZsF69iEXvSc4i/dE69TxGFirnos95aIl/c
OJkAsHKDzOs5FGP1vDlQFlm/jQfTLnaLJhDgB7v/5I24MFVxPNLE2pn+/7AqMefT
V+T38APuL79Pd4cWTwB5sWZHxGdib6ympv1ZpKv1xOo8u52JmH+WSBbTEspUGTeh
wVNObPOKCc8JX4qqqk5fveL2nEldckDE1q2k0/4v7dtPvd7kTy0oJm3ZKdY15Kok
qKAtO34H2iE6hREurWx9gnKao9fiEi9Bl5wbULIYYoCEQxirFhDt0orpsVY3rjTl
x839fH13z87LupY96pPEYSi6beIm4gcL4sC9LxE4eur3AR78EzgRO6DMmvuSXJxK
To+sjh3SB9IDIwpSQUNj4rqvexzgalK4hSSuKtbGzpcs5q//rKOrE0P6ViyQQMpo
2jzH25lPN4pBDnkDq16DmrmJvADNEEjXZ325UisoQfpcT4HByl3oAYw3F80yeIqR
nazhbsNqXHarCXCLBUTk5Dz4G7ouiBxeotYJOiHGoaYDZUOEdZIeGWskIQUkqVJM
18xZ+uOA4jm0HSurdtVynPB/u/aNmaHscz+tvNFA3oFge/Jg+b5UKP9q9ine6KYI
zfZ5neIJFr0pdpvzEUpRPZai7UczK1dmzVxuc9w8ePULe0MTM964vBtx4dZ9faRP
iboWvEXRf27hyQmt1kMLbEpRirngGv5l1e/b3SmILxYj9DnJ17FWOJYcpa5MKYmz
3sNthqHNTd3Izmgxk7MFqJTAy84WCXRuFevHz/tzFR4w0aRZvIm+9QK3DrBE5nY9
7vnRHbJM4qx8bJziX3l4wU7fLUXn3NoRVR8QknJPi265+BLLyvMoDIXyrmXtmDFE
IekSGyITJZvYn3sDrdU521hlRSrZvJo3bBJgaKeUNLHGn0KsCWbkIVSAh45yl+Vn
M5Wt2OQNeBW5/waug4TzB82DKdIfH5ddYoyqHIXlvl5i0xoMWBxp46CpWn7GXtcn
L/7b5JYctia+35PHHr2/wGCr3UvS7Nh3S4SM7PMHwFD6mZmIVgr7iB8NyA4o8TT1
D8vnuiw7/MbqtnCvodydniSaKSQokUcRIpbw50BaNLbnS0rrt/yh00n48RX1lwD/
mTQ/F9r8x40kfktFebyNYzdsEVPnd2lWndY1wlSz4JPAOBxdOAkTFSPtEmJe+zeb
SWsCSNd40LDJALSrVKqjFrFmoGTmN7EEJWkQErzDB8eMRmVELXpSzgX7LhhqLFVc
5U71dYKdZyxv+5TJXST8zPmqdLEG060G2l6SgBXc5cA5eS5p6uoPX7/GJZyofSA0
EOPG6FPkaucStZFQvdmz9Yi4Q6IYbwEGJcMB90VJcHiO6aCFzUuX9pFpNGEGTdYj
l0RHv7Mwealve5eXAyieTR9roRAk5Pr3tEFxGlqy5CBWOBV+GOMXO8fqgoezZgBy
e4IGNBf+tQI+Og2HFBialFoiaJKR+y2eewunE3/CxDMuVlmqesATOM9/0KOLWQJm
cf1JAbfxiayu6qbCLLxlhIA3f/Gv54WX59ECqNufrc/KPsvAXcvcXhIOfwECSdU2
gAAN3PF8JMayj65Xj1OdG7uszx+GFVZwD0/YsK7qtgURrQWV5X19rrUJE3aPSDIB
4YCbXQNHrf47UGm9OML9XyErXeGud1Ks7xw/nSGdJiCvj4fZfVzjcCX8ZWWljGkz
EbQeBKY2cVgtPN+Epu+MhOagaLgGGl8T/YrrpNSE5O3oGdggRoZE1m3Kmvd/55dW
GQiXZzcIKc28raFbaxZ+uxuRk55XLK98AEzVwSYQyA/bW4KrfTwDDAV6OYGDtMCe
D0QL2VaDbwQtqH1wW9ztNYblJJk6SH6h5bKtZ9JaUOCeevi/3mGsKo6RHWPShLPB
F8FB0O9fd+1ixcxKixNYIQXjWiLYR9uHeRn1bAEK3yvFhdXNC6MAewMEZAcGY/S8
aHkFg35SX+MLfoyLLROlNmmWFPWh2Zh+O/CaHfD3YyA/GuhPPswIaO2JRE+UzH3b
imzBOF9s9SBQdOaLLOqwyLUp+11w0ba05DYKhq+bmza83THKbi99M95qhbwTS/CS
vwcIhPkqR/oefNM85HTnzMR60JsYDlKs6DUJWSLoVNFAztWuh+jakVF9Z3hmO7Ex
HZ37meG/nJlxg8VSwBheVcsGjjb9NgibzYhxQkWCzB245WtV66pUP6+ZJSfMXJge
UGZOHzgZNe8gD8y3UGpu/UcYmcmbWh0nvLdyiL7r7K00c8Pc0QzA5kj/xRs/vUXh
Mmq/vv4v7xiel+87UYKQfNLib7PTxZHsfQoKNkmyL+rqf6onnQXlJEzygAdVueV6
ZwdVzsSs5cf2FWbq8nvPeBjwy3XEND6hX34wy4JouDXH6tJgxOFOUNsPmGf4OFc/
cq1rbIlIdUHG8IFhrDOdjznh8wHG85TsBoTnMgHKixS2nVA4LX9+oz/uUtBfOuIj
u82TDZsf8BZSPif7gi4vxU7DTr5S9EsXv9XNCzyAFeBHyHv4tA5Q+F46sWn1Z2cj
2tpYYbOTR/jm7h+TaYqJfNzaBPV2ZLYGDfPrb9UYdJpXcLHqLP2Oi7o3d/vhaGjA
IVQAHUmKjyW9HexjOK5M/5wNrqHHRPflonRUGjC9U3I81uCJqI6qzAFgwzSljsQR
niUmWWGOeOdyAuPYEB1olQlYrsdyicp/+JEp2fCLEBryXuROngVluaWtXyYNRh/Y
BQ8/1c9M2zdvj1jeDYoWnaMnYsHIyR6TK/qWthVvqVzKh7KNVBymI+tPKd2e4l61
f2SCEVc57Hc0BtYSP77F5/EKalmOCP5H6gbsqXWFXCUlOi1Hle/oMigH700lrdmx
ACoIOn4gVn11skmEynJ1S8E51JO/i2vTEIyoi8Od2krb+3xANggMCcgR0autt9VN
hZK94ckNpiBJdnl4Zfm4D/iHe1g02C7bfyNE86LA4VVO7j4emhThkKwcuPmhltfE
S7e5TR51/ykDq7AMFIkZV1EtQfEnYb/AzlSUOy+gzEfgr1pv1+H3waMGxIID5ItW
F5owsJS/ao6hKsyIYurxrN5pXJfMXGygdGV1T5qQPosvab4I+DIkZViQ2hsaX16X
NOhWIdceJkGwY8c6GYi4JcBi9vaphHiwozi8HgM16hNU3MNNCjZMLvetqhjm3plx
/z0AEoH9lX56JB//0TtODN8mdHmjM0PKx/rMrXkP04JIGlfHjR+PQ1LuWuQ2sipr
jWt8amJgz79uaizcBRHRj76QpmVU7Am1a7OsrkMiw7NfDENUdy7PkrhgCYESqa12
Y0nVb3K1ipN6GBZTjFwOz7a+7dRb+K9wABCXEqM5+tJ21zNT6Dp5jmDugQ9vK1Ry
HrwHwdp4uFodxrLQP7jVuNlytY2Vztpi+UfW1n7lJvirPYa9e2MzPqK/XsU9uiL4
GursB2TnlropedBmM4Rq8gi/dC540i+sWzEmvX6mZmLRvr++GzriXmS5yFG3ko3s
CIfoDYnVrPu/BC575eDk1Up6VsWGKaqJvC4xayif0kcOik8BPb8xNgXMIQpzG3a7
OhLXsQxYvi0an/fzlz3B54F3HaKAx05T1wAwHkAGrKYRI110R6aNzAMMCR2sbuC/
XWflKE2t3/Hp5R7QdVPpYVZIyO6y0hAG6eg1RRazM70MSAV9vTtl9pgndi6dfdbZ
lX5ECPLzPHPcy3C4KrZEyY/2pkZVvPluGAuVCK2LjRpELVvww7NI51lSRhjCIImZ
XVXPz79sAveeXnasayndf0Ylryt1YNRrgpaCXJK8a+aSnoDnklDpCLMdZK3mk5k1
46BBR9XazYOHSUHOndjJ49Hi10TuSawFW5q4AyEmr3qzn4tIMbNFXUP49TXXM7EB
GVUdFbboiSp9DhAyd/U30LE/sh8GA99MxzrdWBX53RAtFgnvE0rTH891uA2puLNL
QHC7dMee6GzcGmEje4llzIyu6mTLAE4kk3eU/4WQB+DERxV51aCQNN4sxUj4Oser
aFOxDHql92OCtUtZP/F8URx3gAjYV8DHI577Y6B+TfeGhmWiJGZUrZPwdMBRnuVl
xQ3ZWPBj5FuXlBsuxav8O6/ZfMfTxV/ZJI7rKYQBLKvHHgNFFHSzGazMPm3cBPIE
L/1oJNGgET/utZS11bexOkP/0yZOjO7cygKZwtXYXv1wsjjE0PbERtiwTHS20dcz
zTpotZZyvPLcM9J2OR7W5vxmkEKUlQ5ONuRTeJ6ipBRBzhYqT9a0UQpmjrKXDaX1
J1SgibiZTrER4NTJPGE7klwnF3pUBRzg5yhx2nEz/8ysOC5Gd9kur7whtI0BSG75
LbeFaW2sI5Ob5DyqJlX9UtjuztGCxw7LKj1mFSa06sxvMuV1pue7GtjkkwBYA0iy
pxYa2uq9UoaCfFDBAl6QdPEmgFzpWK1Qh8COT57VttvVbgMbRUpYqTneKCcno/X1
CroH6sO3RtfITs4pZ/mXmbNmZMTTFm/AactHu7atmQ6q/ib4Hd+ESuMXoB3GvaiC
8YO/xSCJBASu8H3Eq8F54WJw3r3rLW8aJVB/oBfPz++N8UmnoPpbEG1vWXyvbcTQ
yjFqPrczcb3ltA7TGfPxbRI92o7yrROokPdO4sHd/DzJn4i2ba+tl2sq+nIza0Nd
hfDbU+Q34krW7QEphdaQiyEf2arixTgs9XCYpWcBOEtvWlgR8RtIKAaWwu0htpPd
LHdrAElzdjUw2OL/p9wU1K7ug2ZmAJSm4vQ4fV30zUYIbQpxXHlMkt6WszKHLM+R
L2KzFxtBUv6K++/K6RghyO2fkvns6tRCnTP2+iv0yMYNh6CLq0f2wRsNMRg2fYkM
Hcn4edrELd1rktzVz3K37ZKsf8dE9/jx9mra0RVRuoqktj8lVs9vw8WKXU5irZOy
zblE1IC/kWqPLmqnfUhuCySmHzDyIV7uJGQ9vV4SMr7bMSVKMMe/DA90HZX+oclj
O8VVkPLlun1psXo4vjdHN7lRzBN+d/KA6Heex+CPFADoN+QUlmRT9GzuvYVdvXwo
K5fD9n4n8FmR4mroEuV9OcRb4UyUWMUTvDu0P1n6qfQ12j50uqhrMvh/9IFJoLSW
lyhmjswdmt3Wfne5TqXWzjdMTai4uMgECdtg7UYsbGTY2yAtmZNkLRNhNffVSoVW
QmqKJ/Fb+VVuGG+0kf2csZFFWysOZRhWTqo/UR+JuSn9RO0b/uisNuqfIf5tNAAT
jYvxui98/NpWvNvlHtsSj2DisqPRG8ZPsvx19Ib1lQTaQzYCtqkA7k72SP+6AbGs
dVB2Q3S3lRgWwFhEmzTb80J+qj6d3n+0GjJM+3EVp16Jx11z+Ze1iPcgL3KGvMbm
cs2OeRjd7sslq4u7/5XdJSse24Kx6I41CaMD0IeRrJusQ3bwJjxRcB3DuNAcNERn
QlcgQwVENelC978UEqr4AM5JvOd7VXVGqxemlT3eohvOqFEjsngc4OKXUui1QlSz
Y6VZzynUGA06D7BAJck7inAQd4LmuBfjLQ6NnfaB8lSYIfiNu3g2cagElvGMJ38e
azjdwu/uFsuFLzKKjzZ7zXkA+qOicQy7uj2FNUlyjlodBTE1vWYBzBHrHN/lD9bk
7JAqBjez3JB/DS+LsA7h7FCLkNsGHdD6EVIxDAveh3bmj17wFo8bhWl2mp7cjVH0
xLEKr3KDek0nn7sa/2Pzg73AVV+o9ZjXo8KSiUOVcHQIbAYUFKfPTNK0H7fKce2m
bGQyb/OoxhnYd49abjIBTlzL4m4xZJKuuQg0rqghrqOIi4LQoFuvQKZsF+mHVT+m
RbKdmN7EaaDJS7RWnKXvKBMWv8ZRvy+c5BCuBt1tDLANTzWxi0fGhnOOWirQBd2O
+IBjzJ59nvDRAVH9nQwx4XfuE0T7u85v/JLJpB/pZ06ifiWoKNyqKYQeBgNN9xen
RXv81A0sHoEJfIQSfOwk3NoTMSEajLlmEjY+yWz2UM/F02GX+aRnCsnTW4QKK06N
D6pR+7BCNjyJccQ3+iZ2PKy7LqvkKWD/BFWYAUHpprpL/2MIN5MMLp4tyGfTFdbz
EubuBLvyhIbjwLn8uNAmtkS2TOzh2whCrMOTwXs71Z1iJni9dsz2oF99F63h979r
/rZ8KXo+mXyc4r9urdhithsXhT9DMSF2PLH+soWFvsj+E3L9cpnCMz1eZRRL0Cwp
Z9W6EZWawqlAECCJkQmHZE8ZPURs3+NRRPGmTvVflMw0oXBPtHhuNzSVCMCs07XV
yR/iAZHajAqaA2URx0PyRdR8MMQR+qpY9f34J+5sj61lv4tcx9ZFYP+BfUm3H1Xi
QFz+pfYsUFlAVVakHVgUTdBI5wpzmXbt7X+NqV1+MiMxIwoheU/X0QZ1ls8uxOjV
7BAGAht7MffRTbEncPSE0LiNzB1rE4sHPl1hR5of8nfhKWCCKctv0PhPXicQ02vr
nDzhZjiHKponSNh4r4bsa4ZfTNwZQVLS8AeEt1PrMhgUMPRFD2m3X3NnLw2XpReL
6YulwSYeLBhne6PC5fKnDigTKEVN3OklLqooqvO77uXooVKz3i0IsZ2OGUKK6NYG
rrJXcKBW1ErAl3oI9D30Rw65xj4d87MjoVwX+bfPKY+/h1ArQSvLMTQZlR/pBNQa
tOzJ1O7Apqwth1LXKJT39kxHznC2t1CiFvGgf0lgnl1jCky/Q0Dlv7xJk94VT/de
PaHgud7Sx0Nw5Nu4faFWJ/ayEig3RyMHLyXe1HPhgfatpkhbmxz/ar754SdgJZqb
Qu5AlcPgGonFv5dljE3+aCVnaAH6i/xJH8bPDJZObcFuE7s8O98KtSSibNG9RGow
AdawCmNEB1Chm8GYQmP358H2tFk2pKiIjSGnBeiF8HSr9/nTkSChZHVzC07ItrBf
E7QVx1d0XadJb72L6VWAepnP+FqC82UG6Calx/HHzXKvAQtAMOI4mx68hb+QuMIj
LvdUQPEnEN3scgD7fiYPOuUltY67JwnD9n3LnqAfzfT8r4NPmbLgk8EfBvzPYoqH
fUWnQ7TF/7tf1HqOAoHg/Ft3zwZgvtu23UlaFgBfzWl4lTA7UJm0PL3osrUWT1yF
XRmgmMak5uKEkPQHas3nh2t7muX0rjE5sek1yzn+IBKNkvVGPEZlheWJUE69QdwF
YFGDQitezQHeUhZra0jbdvMmALDo1ggM4jIdsWd9JDdDd0/JbKDpujTflgU6m28+
P+xtZR0RHfWwGjOjrlv5YDjJczR9DCtVsc6/WNNrqUAP0NB1JPhpk6+pQt6roThk
L1S2xF2TU9fBkdc1mY74s9tIVECwcLXskWOCz3xBHni3AhOpzo0Ugg0t0x+eN///
MZ8jps2kj3xrB6QoUdbGssGywZOiVJyxWLdKfKryaM5K3W/pUNxpdm8beDkjUlrx
DL5eTjPsF9yV1PH7MwCeMCchHir0tg5BUMdlScn0HvZuojfH+WZEm+0AnDOkYEB0
bSKp89xqb4Dz0cLerFPr8coe8+eMhKrORcoTNdoC4loz3eX6idc1GMKbGZ1eQaU5
mc30jhTExayfvVvVjWZVHG24XSd7KFhsAcaSrEnN3K4IONxMMW7nqrf2EvbSXJce
oBTwwKOpm1jukUhKjrSgyeOoJ/IUWXRjskxCygOmjhYQzTuQClYXaT5+ERa8ummJ
tDi/EMtRmSkM6r4NBV6kb+UIBE/oHmv89KKbzIun1XVq5ujocaVLEqGcb3JJ8ANP
Ufm5cxzjwgdqIlhLykZg2lz/E1rBe9IYeH49da66dpNz8zV/43FvfwjtJ31mGeuT
otaMxpFomaab11UHtC7BkW44zlCcQJBaIML3/amfvrNE3mX2Ju6Mw3MQ7sVXl2kp
c8wXkdebMiAMfit1flekO8fo+IVLqSEXGH5O8Gh6w0t6I1eTL209INyNtGxOLVmr
dytwih0OlkXFO+vSyhWSHFXMa5FAUhh3ACimE/XaHi1i9nYVe/kE8ceyV3KdYZBx
yNFgZTWuNaJqaMKHSxhv9RpkZytu4fR8jdMvJ1vTjgTQPG90qBGV18c0tI6pzdam
TkPHsuUMSuUojyDiFLJcpD0+Zv/mlQnUGiG2sGaa75jAPLjWwv8kHaR6vyr3B4sA
2pjsomgVOdgfj/Vg6higNKxQvmMLQ9Re3+BnYDjDlnn3/Eqp8ENF6vsTzbEM5QIK
yYzOmCQGcD8FNztbJkIkyKohjZu8rUlDu7XibnpMdV5su2+/nOD2AW6FSy01YYfK
jDDY5UItb/RlydtO4iX/kOtyevfjjRERROYYvWAny4Xi8+EhmFlu6wEDZqFm+xnt
PHJnUjI7jH10wzQ3i4eKW1FpivGA4qAnE29IsHurtyF0fZra3V5Sxr3fc+U6rfmQ
FGeFhazvUuLzky5m14cB4SJx2ioaszqzIVmrUBO9iDFHPed1GZStBuBVZAg9+dSu
DOqBmd/ZO12cpdbYPDhtv4rMst7PhPtVEm1humFRGf1zO7fEbG+JBfvg0xeu6kU2
pGqilS4S+FIjbT6MuG3gqyTfyVRJF9BdMBQEjbkILf7TnX0sb6vb0xNIvBZMGvUa
PPbLGMXjAcDGejLDEU8Sj5lfVjovMELRTC2aHiTk5x337hJvVstqnKQ1eBUy/V9k
7YlqSdfARKmGCpJvcwBpgvomANkwrP9YEDT2FxSCwzJ2E8xBNSr+hnADv+05oYej
rp5UhD83p9c60xqxOjzglFLaXECLTZvFnVKNkcdBKfrn8ALOv7ZVcKeF6GBM6Ujv
QOiFuzPXP8nUkUaRtN1D0IPi6DNzrq6F3XhZVxwtdOeApOvxblO2SnBJeACN7OuG
ixZ9XpWzazQhDwk6G+aRdT+WK61PXQZ6pUlNiJ/4KFN6edxiVDMOuyq/WDYvIt1c
pR3d6pMHaj0N75LxCd9M/9XsKJ5X8YJtePNN3IXxQE0jyRAMweUaBKBRzJONwn70
F0eKyG2iT6aSEbpGPhwuwOvXWAsF0167SYFwLFuO2l2/9AwlyjD0b1x59LZPHBMH
m0lidR1SYcRIsSCeLBlpajyEW/5+9ES8ItCs5MyjnIxjyl7PB5firX9l6f5DQEsg
FWNHgD/6dmdz12Pmsq01/d7B+UR0EbgIYsmVuhUFTRtEA1iaTRjQs8MOMCK09ebf
sPsCG6jqPIFE6DjS4emt7PLBQrtGd/ZCQ0sg0SjlrZE1qOyoBlIJbbUHWLlic8v7
QHL4qKBlg8biP1xQkngfIGfdva7K//mWnNM2p2OI8uNfV2YNUIyRWjgnaaIORgeO
39W2FvMRSY70iPamvYHr+IRHywAeS+FDLAJL9HSWgtB/+3SkLIXH3cuRMTlhKbHD
HnT7cIyib7zXSVvUD9VqmWRxo5+C+WKP7vjkMkjcydZpd0XChkRvZnk8dQJRX2Cl
ymLMg4qMUoQeed5yIpzDYzdRT3LvJJ5RMiHmnFidwNxiyK0m9CK4+iKAgLel1JWp
gs+0ynB+K6VQPYQ1Wdph/JFs/VaRjILr5nHaHHxzaNy+zEJiXtbe2WC9yEB/gOHE
SENfZ6Ac+TOiNHNTbHfEchhj2dCpTuTu9hbxqfqbqHRmfLrBfI2PhtFO3ISsPZ8I
ewd96Eym+vzgy59kCJ7UFgPBOSloMHZ4R5UlOO5r6IJy1cnhWSDn7kwPTh68L+yH
lm0n55vM/IrqK8GUyUMhY0x8rNJ7eVHghj3wmwkLvNDTfacrMDOQL0TTBN/jmCgk
b8epUxdRB9IC5bSXX0K509IFY71nGgS5DqgKetzr/4nwCs+DoQatNAnR3H0f05S3
ymJiQYM7g07DrhMmLmz2/Bfn9XwlDCqfIvJCalsVp5KpIiy68Nua5bKqhb29+49j
RHb1crhaZtQMpYIFsEoU2NMn7NrDtTvHn7XFdKhqIc1/sy+QoHeJoRkE6u31FDcC
05hPk3BrSi6IZZQ2/G2iRxcI09wB5vWcQek6Rg6ckDLFEGLDpMbEgoAi9oNKeYGe
Ykn7cLkJ2x442+HkS7UFPNul/j6mCKMxCvWj075x4YVZ872qnvMKGpabH4YhuZym
wJ12JaqZeiKLCQPsJ8gPDxHY3ZmRtonarK3ilLz3Syh1eXvghIKfUeZa/9YUGAP7
GLIykFPI7P2yS59tfixGhypGHuZXgAZ8+PhHwxuYYYut/pBQ7rIUlUZwvp8Tfkbv
BXmTmKs0lQ49y/Tyfz6nE4qVzdjb3h1w6f0BtUc3L55F3kPpWAAoolTal86fuwSy
DdZJMJrhPvups7CI1VlF5q/0WCbKrE92D+75C6l+7ZCh7/+Xai+HO3psxTnxuvSN
hKk+BtS0fFF7X1pBn8xLxwvjc6HNm+C6AekS2oNCe7gadKlB0jZywsc0qXNP/aY8
eG/eJ1S+Xi0iMPuGlS6rQRHIkhqf/Ryi2yWjhb8PLr7IjvjAxXok4RJY1LtCSwdr
ewtr9vLCSv8nW/cJFBehix4Jm8PKK7YE1bKiwE7ztm+46IkQpUnGWidRWj0KLCdE
r3iRLvOVzeIJE/y/6NWzVk52sTkEkuIz4cUYg0lXv/b9jOpNsEgp9JSz6VRV/Jde
DfOFxbjjWwV3TYeqUirySkNJGnMa4Bk9GF5S3TRUW4+/ntIQxN/8C2u2Q6JKd86b
Yfjn9o5Dlrg7onFgSNpo8cpOfjSH/ACOg6elocaYjtN0atgySgO4nH1w7/C9PgRM
FeG8zKDAaLUy7VWePlfi2ir4o64drkFI093hq1Ysf0S2TI/DjxkJ9SjiYjOXRzNg
iM+Tg9mRQZBLnl49rcne+vHFo464FgFHo7p36RPS0n9GKIHnxH2X7yT3s4Ky8ENJ
vLyPw1WOmW6tXm/sZ/Ufi9ODdPZJw2zPyK0ihlf/Ob8yb0mE3RBVb7YAxH+SIfYf
U0tILvO5DmZWuz8JDf4LqAdOYKHSJlPtb1jMvkxmLiqPs8vNSoggastR42mi1+0W
uY431yS/UQs+8bcKwrDXiRd8HqbknNKBzf9PQJTeOIdMljWqoxg0rvG3jxV5DOPH
z8S3g+8kVuDG5oiQwbbQr+xtcoYyowheOzQVI8FdZNbEQMMX/8XzjZRhpcQPhKhU
BDY51Q+PAaQCSjhPBJW7AkkQmHuA7t1MotKAcW3Npx70vRNBVwuCzerI8kdENGM2
AvVH2gO+GRPmrk1T9O+mjACqiqzBtVxITPyLeO2KZ8JWbRa8WeH2uMvlCFnNspCr
3kZdkKvNKp6n9Ozo+iGjFGBu03S45PpwOjJ+JigA+o964ER+SoHEvYP/PmyYjoLY
7msVppeMyh1h9kM2ZHLuXZDq55Xgyd1Dtnsh9VMdEisl11Wm63KpijidAC6JlQ/D
wpGHxV7V7sgcMB7i5IziyUpF2EWXORLwRgDsDTLURILwWp7XIO5/1lgSegizbW9N
UITCkYC56gjEi5WUYmK0RFDyy++EJZYc3mGhFJ9fbt421RLbw6bLSbw7QAwrIljV
EN0uW12r3IIFBykZLyHKy9lbyCLwVTZyT+1tflQOmVh/Ae/T5ryFFdRbxDOnI/4g
4WVsXPdvq4++soanGWVYhWk2jO++IFVgR9QU2x957XSH5hFL/IBw4qf5qiEk9F5p
dC3IuTAT8Cndn1aOKiB6/DFCqnf7C4XPBKFQA0nFsHaWzNZ7GxpTwAIoBm57Q4ze
Ku/Ku1NSmoL8dNNnKB60r53iYf3tkp3uyUCqkfydMOKSJzb4OZuxePS/ijgLAjC5
b2BXvA57yPwVMtJbotjVmRyc/6/qar6CXsjdNcEbv/pGPqYWy4faZVxPfqRMk1Jm
JjeYQ0Abbyd617mlEJu1ommkfi5Y7lrtD5ziYO037EabNjNOq7idzku5T2rukkLF
8KagGc6+aDJ6SeIFtMoxkIsJTee1kq5M61GDoFeA2VdOego6eZ0wxVx4RRoz/0hC
kOw23fmNjXP0FQcNxVbXUS/bkZxnQ1hijWr3SZJiR0z5/2a9vwHiecW716hEHAE8
Zg8UZuOj9vWOeus/K254NieHnXGKi7ccmobM2DWSjXDvJF9NKbBczkZKW1tAhkJ3
zLnzoqPQn2m9MKyG6DsBWkBrKdJ2mwgm+oMmliofZiesbPIHk0iJHnZzW25U8FcJ
jKqecTw5idG0i+rRePX2piCymi1/jbAYZjDjydQj/z/7PQKwplVkaWMPjxaVfR8x
G1b4RFoOBHwfgCSI27LH6SsQjYIfcKWqeNRx09gKLSxQ8ztQNTFPjThAR9bsfaK2
Dxc6rx32L+xMJ/vAxD+jEfY2tPYsthIlScMbBzTcsDO5Jki+kU2zXhz8tWf2E+ry
o6rDoHIcTNv3AA3WWYEneEMfZ/JZsWkzRwFBMZmGHoD+VapFS+Xj/gZZq840xs30
yCr/sY9PaDSurK02mKYWLuOmPDvcwuih6t1QzbSUxoaTl2BCnhth4FZdcfJdESaw
C3XiqWgoTWfuIx26ImjCzYTobBl+SPxZhvTRG7cMCps+GgSVloh9kPBAJZK3JZz7
Tozbh5GoRGwyaHcnacm1QWJrJsxHytJRU14dx0J7kp2X3yEoxC3XrRNDKwApLCYA
6Hr2zjhYupRz3k8QkPdOjbOsSWivUQA1rkd0yLxmC15kAOCFjiXv/J4mXS3Pej7n
G5ubRtnecpDKil1L90NWjcGXr+r/Nxs7Mw5niqjV+LvbouP0qRECrZ+LHtpK7Vqk
64woe5ImzmRGLq8GvHk9ctujxZOFoMcC9RImLS2GwfTGyMSTKy7zwK+/wqam/uE2
ZIABII/C9gAXVpUR5uraIyCSvNR1fvTkPt+5Eii77+UCdeVJOwgoFCJ3pn3x63p+
N21pwC8XO1Xtrjj7B2MQuP/fxNrDit39x3UGbjb0HzbotUBKIwvotpXSWQePKeyt
gdVoWuJ1rX/CT6DS2GaIpxsIYzI1Rg1gJ/dhC6l22NJVZOpJAIY4oTAUBWovgWgl
7VfUHnVXP9/gXaxZ5n+KScJm239OUIMui1KpEeWK5AvSESZGllMqR0Kvd53Nttd9
9SQdsEhIgFOpi9aweaBK43weHw6oJnT4zSxY5wINLEAzteDzi+1sVDIsPA5ScVNo
xRFvk77I490JkE8zo9Hc8ougX4oaixloch84ERTDJaVvF3wvrtXr4B9DHSUNl/ZL
djlJDK9+1JKzAHpYwU4kdy90Zga9X3Z+FCe+7KvFig4YDIAhmIx4uAvfT3QlX8Fb
F6ooYd18glofy/Azp5Tfpm2Mp80GlB3t0OOQSFxctsswRsrU/s2YNuSxQCKtIiZa
uI/Y86MHXfzEYED0Q9B4mYcYZ7hTGDtf6fVkEhfG4OOZARCGTeNj3AAMf9+Kxxkr
npse6nAxOZDozKsy+RYMtpdAZjzCY8gjRBZtK80EDyGA5iTqffutNlRr11s8S6Z9
r9JtEzICRQo1a9TMFl0IqB3eMjUz4W7m6bMTE19Ph+6nGFQU7sYx/BC26fCrL/nr
7d5MUUjePzQ8a8NVXmtgzDN/PQoPG66qtDN5RFdf7RcpojzLJAfQDA51ThE2HDDt
poqAw9h0siESMF+zovnrQAEhXbozr0lZUZJWLTeU0itwMM7clNfJdCGmG3O3ob2S
wgrqHjsIa/4o1Pkmyk30EluUEDA8vQXTtdSc+CzomKYTZitlndTLtmOL3eIEmre+
1CZddui2mMrVtafKCcbmMhqsr3HwtsznH8xSSZ/BYXgpjv6tMMUE15ZTM23iz3F+
PV2YEXUAzltnczAdKU5JQKCAiiFJBZDDzRlDFg1WHPcNdEYAGWr8S0OiQ6pDLw4H
G9GEKp7gLDSXhSRBrQKSTCo4G6yjN4DvoqtVCKaOsZWAqrdRmB3m04hlxQiv+Yu+
x7/8exdRQdghhON2bOfFmx6QDDqlycJT+48TBfvY7Pbf+9goIvJwXnTooRv4na+s
0IKI7FGdgKnr/3T98Kk/W0jHaycEl8Ldzk3sqNiZeSU2lmP+9ToHellK1Qt5waQm
HJffcU5iIgm7qraHD7soMWVzFMZjQSpVpGa5/R7KcGk9AsCGRUT1QfKIZTuPbnHI
q2lA/vUIOQNThsPhS62VdHR1758uQ9Dncj6Nd/kCNLAOQjxfsQ76skZyHMDDM8pX
1wJWtc5RsHtRub5R8qgUmvU2fgIvBeaFTe7fuKuS7YO4guOzyzzz9qv0WH28fFkf
qjqjt1JcHSwS4PgLmvfBZ6haQUK/BW4YzibbNxxzTpSnjXa9sauYnUMqN3HWIGpU
RZKb+uikvHp2I4XyXahN5efWRD6LN++kVBH+Ljmr4ol8/hAwInqQtPQIubYuUR18
SeJdoyzETc/g2SkUB6s2Bwy5wGXeT9ZVPuYj2Yt248Xcb2CyuT/yVNmYcQ5V7vs4
2S6x2nkMQNv7u/uDPBdWfZhfYkvkVgfePaTburKaNjDGXtm+Dzg9Flt5+vCm7NN+
rBp5Id+mT32I88g8dJ0NNS2nm6wtpSvy7LDXcGZgTRB8ZoO4N4oJ6lw+SeHVzFzJ
SjKy59vyGM0V+RSNLsfMYayqJD+LQjWJLCBfkaabrQ5qj/71GoGkg/AdDRzv9vey
8olMRcaoeajghEuUWwnjW6JBg1AtV6vXe2bMfX79IGXXZll+b0vRmmiqPdjgoXZk
zYxApHKU2TzZ1n1FnSGvAwuscjdZRapwVi7PCNvcEmBiLhiRk4J5nGcopzkCIaXM
lMXEDZCkneLOet/TiSeU7QVGmhH/yvleGqhx2ItX94x2oorHuojif2y+LYfUA89a
dqQlgMKIJinROwouvj1i+1V3x4fjll4lQhw+Cnk6BUuJhym4+TyfuSbsBM2s+dis
UOJ2Me/SmOR/B5sXsc1HzymLHerEIirJycCLG+rBNcwrMjih4xl3O7Z1cMtW81F0
iKzJ7KP0A7YuRcCm7AIM4JnlED4U/smlTP85p19DjyjY/OVrZWKs/pAG8/mgY9dD
mCv+lz1qw9HE4pRGu8VbxDIb9dsOOnZkvMblXNRzuFZo6GBltTMgmR5a3+Dfl2+N
cvFI0imc7Hh9Mn4+aoz2O8cbNp49bgkcFA7C/ZqRENnK2l2ikCut0qCcxhOrTVef
+j3OXpDeD2EsjzswPWuYlNjFk83qM/7tjtkC6i57/8I/spQNkGhLIlI+WMVVARGd
qMXNYMDSX0jSFMv3S8MmVo+Wjn3Ww54dKi2/sD3JyAhrZJHPfDqD8eo4T5dOe2xd
V98IfAmQ2/+pS+1QZU7piO9C9sWX+R3rrVdN+pl0hZBAFad4HEAK3+gxnCgzxxnV
MMP8R6s5OrOVcSEKWEB3DyBowayUOZ6764yLzSyDudobqMmbohULsx+O3wQlXOP1
jcyDgxPI+9OYJShVde4nj9AvCK0YANXVIvNgmollCcNDfH8fzFxT7GRcCPGpicPh
rEpQezLGXmrT/k2MZkIX9coeFHEaGPt4WUsdK261hZlE1u89YWLvi7DcjThmUAJg
e877YrFpeI5+1joReWtV1nRorClBNc+MywTzKGWx6+t8o+UOanJLmUxKK8VYoNmt
RT9pqJlXpYzbRKWYqHXhqnJInAhYtEf2AWP7eu4kNIFc+lLqSWMzfkt2pyto1Pcv
3JKyz/zLQRVYqCXAU4aA7IOUtOjOtnYxhbcFqzwoUZPLjTFmJ5/mqrtVopHMX2Ez
84GhGd3AOssAoDfkVh5H7dv23nh2JHhSNXqpY6Daw/Bqk7gwuWyalySAsYUR2H31
kxnIwp+EZX0hP+2bKA49JL1WdgdRp/nkueZ/SGL0MEOgGszHINnwWanmM1B/H9E0
Bh/aDHKQlP113+uuSK+zkOcgeFJwrKW8eD6hLQEdtbsy47Tn7GwZdRrI6FtmO07+
q3fRnYmR/t5dxDtoTYosCHqsHpoS/0hVQmhw2M2wpsow8SZLxf1XK1HPmxGIhvE/
1A9XrI8b2u/U/sbe1KoUZxfBz5oRZIbgdnn89oXztXRdEwLIUuB8+sWLUeSavLzP
zw0N3qLA0m6S4Kwhezv/EymtlPwFED+fWI80PGVFb0ZE/z6AGHNdcW5B3ym7CUeR
t/cn1CTLtGMWyRTBpmIBVcl/HhujlX079dhAVptDnbJrGMo8OxKvQSEIvx2GTW66
JhiJjtueeoBy9nM26BkCTprw7aE2CNlbuCf786l+JOB8ltczLBnSzDK8ikQ6tCJP
CEiouyV7ElGSiNa5pDtOK6+evphd4Z1nIuQ5HmYN6dn7Upj3M/ohQ6zvrY+LeV9y
4TiFNOQ7DBl8Pdr2ptHEacnUkEzB3VEmR0H5ZEffVlDmcqP9b9HmQiO3DMVFQVVw
ATjk96vhdSzo3LYlAsgfhNDQxVoUkypQqicPrpizixW896qk/pjfe3rMelxXQtPE
NYdUGiJvQpR1W8S9ziGlb+JEyuiTxEzq95Y5rxnLIVDdR/gCPdYjz3wfBPM51jm7
/IUGxNiNU/86QCagMjtW5Ui0H0HIxdl7moq202YqvSFVYq4AaHgcDipDn74+wJEF
RKiStQlVUQlbQfODLgYV3mfQi/EYISaQxiOGXhH4f68znET6t4ODIMyLBAs4V2HP
uF0I96quoSf116Yb6yk/O/Wo2xZsODW/bHZDuVib5bZyaxESwsg0hlUndUFDpy50
h0V9RTwrAlAnJKY5JUfCNEC+X1KpK8+tlX7+6JtHq91IqjrGT8pPk2Za2YKfdPYC
RkyhjM3A5/CcXuLy79plXb2iaOfpClY5E6YCmCGnd67GocKtB/A0iOm7ExYVnwNx
6tybMuU+Fywzdr4+hB+WhgaCkTwJElqNJ60AcYFxvZWwVbxqmoPuI6nQzBzns40o
5dtTeSTid5FmN+RznOIVyUD2w/bmacWYks4y6taYo2HiSRDfdsex7oEnsdRttARE
GtwPb2g4lbJ+TW7q7KNGf1xChviG2OuNATS/XQxpPAymSTxK5cl8w9PeenGEAH0P
vDp84DDBCJ+D8GzT8YYAwzjBSSDu/HnVNQRFxUioQr/ubyXEzFVEJyS2qJvqNgyD
2Bb/e/md5PBSqpw356XCGBM9r5ZsEjmqhM+/LWo7IhBfSSw49Xe1Tx6GuIAr/s7i
taAXae9G/XZyIdJ5MpTC0GF0yeVY6d89RafqDAA4QdQWnh7oZFZvnxW0wg/R85xI
rG9c389JTk3K7181J4jbKOvlg0Oos7zuvm540gB1vSZqr9rG6uY1WE45TOfMg0A0
LlEG6iCEySNRIx2yjFiSK1Jcj5l/4Tl9dDjQh8rlD1kkDof5vIHUWmQ+xYSabvNC
iJMVoxewfVewMbkGVD+/u8n5mvUD+zwXagyFPWyn+h8Qkq2rDZ82NTJYNExatJcT
BGcAvcgvxKTfDL1G6H1bUILmZD2TekudztgIMWCaDPHLmFfM/8q8wEnjIiKBiDmE
CK/ryiTHYC50M6Mq1pfFGQ3mKW4spwmKDnVqMSJ6qpxFsoga5NtmCWHug8pG30aB
aUXIIw9Em7109m9BruW70lyv/GCsALa+VoXYtL3GRlRV/PYohiZeEci8HzGJFJTU
TmhBDC/P4MZh5bwrZjwTQjvD//DwXxUmhJ1ybu4z3Hpgd4ooUO/SLByAhSyP42Ih
UEAUcE/Vv6fNBz5ArLMtp8eD9vjiz9CoqNiftSRUbYBREgNj5bG2yZrfKGUWlFfw
/s/zqh96thOVq0bvs7YQFUnEMiAT8+o2xVr4moYHpzXlDScujRRT2ylz76gstHGu
Cz9HenJYDR8cp59OUmf1v3+hAhS0tVXyd2ZyrWJ3jpKaTYc/YqEYQmq3U+WkxKsx
9QT0f17GrODSaSux7bPp13i1lkKZ6i7EJJCEznupR2S7Y5PgFUEfklkwf9AgSZL+
DjIuRDU1CLXXt/7CGlHeEf0EQj4oouE+trzkZcJ8DkOhnE7/CScTPaIifvwwk7fR
hCJO0spereBs8ikilafqE6s3gvw9usojnJmE8OerdsoHvQqKdRkNet/V8DaPiwgL
FAF9RSVwVj/+26e3KKChGkNS3glywntA7l5AfDx+59hQAKeq0/yNtK0PxLTq5wpM
5DPTbByUr7knxHqZWEwRyGo3jBBJEnZPJk2R4+1pzqSWcdkJNziiLL1GwJEU5YNg
A8fT31edYnTZ42cK9PXXH8FL6I2mf1KS1PZuM1RRkAK2gaIdsDIwCOz6s5DiQE96
YHnmAl8Yncl9o786kWfMijIlitABfDvi7oijCrnBdvwFHXDCy+trGTPpyCGXSuGw
Nm3lQv1FgsFP9Z+k4Nc2BVtvjRsDYSGX6W0OTulkdB347+jB8zX2zqoMVbNXFOXL
Mg5nd4mcWTtOotsgYL1mG1uv1XXN7XO8vCJ0pH+bKAvdJiF5zKJIqjyJ70gaI5yX
7F0Bb01+7G4jyB8i5otycGZ36osZWfkWo0L0F8YlbzeHQfuWxaBrbmXYtXOUJd8f
ylKMsvRqiEzOkDrLm/zxHGILktkdhvxNHMi308VSj8MyutdghBEE+9RfZ6UEZXVr
G0axhg+F8+ySDn56XJC6Wac3GKmKdjOiPUlewSvEKChj2OFVvnOoh49f/t7eCC3N
VeJlYfugzwozTgOJK1fIzWN8uZLMYw0KIoV7zGZ1FBYit1p7PKmiL2J1BaZGnKPE
Z2QTIsGOR+yn0qNc/YRMZmA+Z/irguugyvCWN9+smxgjYhy+0tuNnxw3RitHTp6l
A8hdJApe/mr8TiBabkcLIsJ5lMIRMFXEkzevBjd0DH8Ux8wSlQHEUWbL+IL+DisU
EWhw+NBkNrkrpqKXCF3BD+lAwBDYEYy+VwrPoDJpQEUGkTbs7ux4g1BSUNd12pkw
Tw31zxx6G68mszNN6iJ4Zyr6YeoduvBNKH4HRtDXUThcSAdDErAzi86t9TiJXPOe
KMkp6F0nTusCFR3o295Mnqqf92lZT3woNdpmfZDA2aEbLQeKMi97g0CjHjuGlB7f
9p1SrbpmeF5G8GXBYx9tVTm6ViuK7EUl9vVOtV2iokJdpRdZsxW2PhvjT49PxXZg
VL8d7K72r5V+nr9oaLZv1xmJ+h8qVU73Nw2sYHyOAMwceDrPWb0zs8tgYKI23wgd
Q/U3EwyPnd2c1hSCySQhevlOCX3IfDHcW711ZU+wgctF7zaCF0E/G9jJnSD/NYn2
z94dz9DHIHzOXwnkrM+qJjuEl4VzDCmRrSENOPXo0YacdZ6MpYbfpo+KCH0kJSeF
4T0KrLvTgpXPwxXwYBlw+gYsrZTvn/to8bGDLB9iSptoSxeP2gL3pBLH+wMvIeJ3
MtEonwzniW1IaLHuJJFesZ0Wigx7PE3cyZLa5xoKZNrc2GrSfgH1qkPE9Ke+TD7+
g5XWccJrlL5RYCEUGtw53VYMMbYkMH8vmpyVKYIpzs5shErk+Rx0/olZlAfUJ7Ql
TR5fj6WNMzzQDY2hByinNu8tP7weKQ1yrW9uN8HldHkgwqNUqiISSKWt/uyXLeXQ
sN2owl2mLCtDFjFzeViPGXOEo855FTqk/kPBry9WW/mWIZ0nll4PvR72nBPom4kv
DKgo5VRTUn8rHnAFLDCtUH9hDyU9RjPGCa6oVI7VgYwMQljEli2wyKAqB977FXHx
WU+8UzW71pQUxSGmcPWhO53AXiCdI2i7/Nl13J61tDpMM54eH6epqaS1Tnm4bgQi
6usFg9XpcogBJo4/1SI8/zSIbB3Lox1QxjCrEzO4s6EkU0/JIG38PmQHLLBDrp8s
cipJBGI9gmCZ2WeuqAHdDoMuKtmQTKYp0nyLthpar7achgHsf3HwkiHbGIWkUxKA
uj87GzCBAkfOgVz6IXAUeiI13mIFA4OvLcOgVr/6v0Cpak5xc3sWpZK71FzK9o+n
GnH2XvPMvUPxNGxq7u8N66l5JZMYMnbOoz+IXxTxoBxJ3IwrQ0Y6sJKAgE1qaOWh
Lz+WmUvhM2V4OlHJBdIpJJAV4s5r6tsH6yDLt+FtxzsJJhwL8PKzfwiXMKOQ10kO
tp6ba5tSD6LTF/ge2dDCQVIm9OvS/vm/ypuQVnrRv2TxmgqxJo31OyQosA2SDG+C
9TCWRCAOf7+FPc2AgiPoUCthwxqkdDLMsvFm03H2uYl3VNOJAQozhs+au+HxqCWA
OWJldw7ePaZ/iGMUbjH3p74mKJG+PR0LUv39q1X8IRHgYhTGUtmGfO/7OB1ql6O1
4laLQVpG1z6fLMbD7g/fEXQD6xyzJkxO7QWX2PLxbzsC+PXpk/nWpCekir/N6/lX
mZx2xSoSKy1DpbLahDgDK+uvF8o7RvIf5BSIWiq0n9gWECmb6jpWH4u9qHcJkXRO
U7VODqaYA5LNvY50s290z5ZZety9WWM3cYirQyh2zIIOlKnwpjoqsq2D26aORvG4
geYAozFm/I9oAYRHja8UdCRcSgxo/mgR31xhpLpc2McVKP1iMlZQfbcnUy6sYvyu
dvk4f+z1ouxrXOBA9BrAxkcWFTkTOqZGHMlr6N7CesoZxnOgGv3ZRffEeI2g4IZ4
k1d+F74bMIQs398NnOVHr3UIxq+ydE57WOolwxb7ilHgCfkcef7dp2aiN+FyxNvH
VXpZ8QTC3gSpQH6y3CYCyOJud3UFDghF20xzjUslqjke2shi0INUhfDuquHtdQo0
MQ13PppfY/EGDyQOCvPUSyLxh5raITECjzx9FTFoywfthrZU65ux2iGwS7mw7hq8
wpWeHjMN1Pj6NCIyxvGlWqSe4IZcXJcaCaYW1ANfCUnC3LNxOxZmkyGkK0LFPZ+y
5aHfDVOAqRtQjMpDShHdbbRjj58BLA/NjWqH/sD4OheI/f0k3+qybbY2MchUbicT
VYpGGAyv6BFolKRfgq3fljTsf4XnB5Gd1D8cIkMNsDGfjE1Lj6rtCrojHVJOCP2A
bbBWciGcaki7UyfllLcfW5Imhk8IGebH16Odx/VStQaylGRLXKrbiqQBpyFq/Sid
D0+PxXfxJj+0i6vcYh1IYTNfp2GzQqC235YJdeCJ6a5s1SpbDYVvsPnyPcCWoHOv
q7j6Kl/O3XyAxR6oAlVvAKTBDy+u3zbapfy6gAIwZMrwCTapdXH/svnkSCC2r/hy
GK6t0Vg3RSsTXjg3D7Moe+/Iof3wcqWbMdX51HhoHxkGaxjcN9s9mOYnU5LD3G67
ftlZcXN1pw9O26rWCmjrO8T/CiLinFo/nuGp9q4PjvokxAn3Gx78p5S6gCF+96Z/
r0HtyVULMVfCMiJe7MoDPzEGmlfZh7662WM7U8GqJbyY/pukNhuhmUoSl+z4H3Zm
aRmn8WfKJ6ZInahAd40Y/KgDboJQp7xlnu9npKcTUd18mjNyzOTP6wVNmjUg2VaJ
ahWQDUK62IXt/DidILtPK+2EjhnwD49fwvDde7uT5k5fm1KFOKoT3wYzY7GbxKRh
BVZ3i25Unj8t9W6VZBNCc0miTzkCvJDfGo/oZwOCYTyPeKK0a0mFqWo7MChPb2/B
JNVKUNJqwDgs1nlrGzR4CruJwIkltU+sVC7tar/kqSPMcaFCcXO5GpHk820WCkNa
/nJtwedEAP7b1/xP9NdCVLcvHnilQZAxaNlVF9YKd7iFQmLSzY4LuNGKuxvX9s3T
VZwG8a5hNHqqm6DEdUB+d675k4x7BQRaDWPg+a30qEwO4R9TTc0FPOFxRjMsIII2
8QiVH1I3qyakzCgSvqBt0ZGRjQyjbG1C0ZdSbSdupoLCJ3IuGCL5c+r7ovzOTOkw
DKR2yc0b2FgdEF59q4SGx5SsVRnBbS8jvJj8XAe1Z5Fgvt6t6w2eAzzEblHYYqD+
Cz6s9H7UjJaPyhkkK3qhQOmdOKp5NhctJTCVawP6wubK8vp8z74/R7VN1p7qUeZI
40wFRukfF4YXX3JzD69Ic59iGg5BBLK2xa0Q87LfpP9TF1IehvZbp4CDr5pzvd5o
hbbFS0u8uwm6gv4s4vs41IbAH8hUBjatPP7BZlGUcztIL427LwwbGC3MCT1KQ7QX
n9Zp/IEpVZ3hDbOZQ2U50MfoVIuPserN9sZCkUyER5WPmmQYst2OPn1Te5c/w41q
HmoncFYFlz6uTka40v3x1feM929nJ5l+ufIwYrkmL0Xmgtv1uh8QMwLVz+yTnGHr
aE+2uJ/inDVWPhp769jVFG2GjgD9c+fGtjLIfPonqC03+wdqYdbPoHbTGq8/OwGG
eQTzKFr5/Yzwb6EVyUSio0PGryXhS6jqpixmHyWjSLrqyEAILLZC4OUYgF9D/wAR
0I0qv3o1eO8E2lLJcUhElqkCv1E9NneQ7n0jJ3LHk8b36bGG6CN3JDL2obaBVHrx
3vcZ5PIYBB8dsGxUSwYtX4VofxJG6Tdq0qp9R+rBph18Y/qQGAOgXYo72qNSPTfp
we4iXgTDt2eoyBuKwgOLRQycrx9THuoW9q7sVmWWIxflD+KnSM5Sx+KMlAgaoSZ0
vsbdtRfH+3doEIMSmnDOk/2eleL1HVJmffd/HyUJyXeauBULSITVRaOS1Eb6WTOO
tgxtcmb+AUL1tNnvk8LIVgJ39kgtBIEVWemIrRn9GZ7gl1nTx4+CdLeBYKt/tl/L
0u9KL+VO8Na14Q3KPhLRNEOH3j3prMySMRe0LWG+IQTYlsodBvl5t+KInC2FAJP2
e4jQo3G8CYF1zKX3TlTV0s/L0pzZWH5HEU19jQkz5ArsfQZg51GR2y3JQFXNr0N5
7R1r7FgPxj+LNnxcP7QlizOuRbuhOR9f0wCqWANhTyw6haWXuI0QQUsz1bxthfwy
aabzB2R6y/diMdo5Z9J8X5pN0+9blz/oKdbkzl6fyq8XfQdg952w0+wt6FRC4Arr
xG9U+BR5nWuE9Za4t+0fMmHREn5IRTdyHg41YfNkmrOW+LwkYuoygQlzk5yx+oO1
Bsq2cPJgbnGjRqmD1Damzr6CY8zaUNmEaAxMg1dNj5gL6+dSQpAMRP9D4uH9AkEH
orzTz8bAWbKCZU/5n6RKiBc/JSV+tR6Q0LKgvNlZj0kompmx3p7bKFJikudWZp6l
wcQHeBdgkYrifXt5g/LRPFu5gdEqhmsO8XSYesgQto0RMQw/rX7NLoBTv/OtVq4V
G6wXp6e5rOoUWmGZm+I6xmQRP/r0OewgjLx0xQK3lQzS22AXOuj0ZGXO+AtDxqeF
7VhFo47iJPoCsU50HyAZpWnrmQBDE9WM2BAEuWhPAcsqZgLeGVmHcbdso/ypP1g4
k48Yzi7HbnmvGPgp+bmq7ZsvNXB2VK9Hppw7yQpLd+mI4+TmSdpiIjiGdWX1csIB
mR9AkDZZfJUXJmnhmaNDqTrcUuvoFUX3AecQv9FGMkrbxpI3xWWdhJghS2Ad12OQ
3Sj8RLEV+SVLWg5GQiTDoiwSHxRemQXlaOTpLvXv/fcqXoKScNp8UedhNk8EUMee
wwR03t+fQxN8uPdhUqo32zYEm5Es7lJJWdJz5ohI/pnDzsb63I1o2ksF0+d56vwj
U/fxVqzm/iXtEhc5hLjIcGij37Lrw0N0zLi+pD3Ugjc9PMuGFH2vsYLWvl8PBQ5b
IwKaCZnu2quErvz2J3W2bY8lCiE/JR97qi53j5Eo7vHtgoxDovq9RMh3yMc41a/j
8l2/nkhQRn6XXp1Xrj/7CcEUD9jF28JAsZbCDlS8e+3wBCMX4CvpJ4whxhd+WyeQ
acVSuVLx0CHfqQiDnWqtZrcYzfKE7nO+2llGWWBwAJiNJPSpe/VoYX4Os82mLyfQ
z8dWdLP8rSJRMMEGBFN9Si9v4Ff1uDiVPhaCoPKspPZ86XaXyBIZ+E523/JqYQS3
iGl7gyYk0RNl2cI/4eD41DBBHtwUMnAE/MLkBu5ejSMpI1XbtOqGAZwV13DVsiwI
kvgu5tUyBNmx9wYc6TEWROouW8kU48UGBuHGVLaUg/2Ttsjv1xghbqaKn6FHhdY9
6wuACysc1oSf6A7/soeAPLUX+G1sCwpSAy8Pv36IY5v8STzjvUgbUoMBopoN9joV
IV2dHDgom3D4dxu+bQ6+Y4dcnPgaekPNNtYc+v89jQ1wgD/9lH2FcDyhC2XgUD2d
hoXEJYig79lDEnLCtBcyFGcfz6eDqTJUQZI4aAK+51EAdnCrjzx2JttYQm9zBIys
8+NezEAvHPBAAEzYRzyQ0Z9qwxIbXSjUdo1K0qv6JJMMnDdywmCJCoifbvi59Dca
Axm1rAByN5TA/noT0K2+PBpXDvjtqXkfNdl5rsziHpH1gCFCb6LaUaB7T7Qtx5o5
K9fcqiA33SEKdmxWLdCWb8HATyF2EJBoAFrVp/Fh9CDBCaD02MThfFeVF/xTgY6f
xhuP+jRoPKeoHOSdlXRflBjZp+6mAdK91SS/5VCpvxCy3Qt5jFky5oBAeXjg9Thd
OvQ50D04p7Q8AoHBCe/I2Wtfvo46+UpTivvqjk/WbVDP1UDhOZJZzlnLgjp1vCkp
x7pt9ZJYz9ZJxDbC0IbheiUWUCe5HpIN/UHMaJdOFmAlwivDZg5DKDWZUiELFeYV
WCZm/UW0bssJbrK/G9vppx4/ntcaxnmMEAB9KLj8Wm4x6aB194FDX01OuOgE7OQT
VminN8vkLOMhBE0VweXf20+S9DAMEOpzzVNJ5ZlC3bKZAPJUWR7TQLuEQZbtR9Z6
K5QPP7sGGKu5+kteQ10ApktvF9sei5az0sjhdmFNDBevoO2kBf4qaM/HVvXG/A4w
WlDmSF80S4Pvx68KFH/0aRW8wOPZinyNUU9NC71aWtmUqSPqQsZTE+1+i9s7miLv
ioNvE84KPXJh4tTpp0v1KBCpQXaw72t+imcJKvqDRyto851WK2br+E3OewPVAtzZ
RovUdh/gb1u8872hX4A9OU0wmjL+moHXIPVbPiQ/t/UTOrwf+am7crN+dmE+i1Me
Ebxv8IHofdzCmO7FiESnm0XjxAyVKRlSj7TH31c8ZQEQ7pxpOJ0MtfRWDeZdDJ5l
uL2k1fMkF47c8HEKnlJRs9o1Zg/u07MKHbJmDcIoGfwAne4ouo+Vs1iyw+8Nlc1B
qfGPB7pMaD1wBrCkanaIP7BTrJ8KwoWFFGgr43TNwutrG31ciPRzjQbRkku3Ym6s
PMkFissvFagTnQtupL7bBuubq5v4mf5tarQ1t69Hyf5KS8KA2FcozyA1ZBw8FFfd
+ZRWvTeun7nk2WmXlMbAM16dz2ZUJrXA1D09yHYWAjwWj169d58hd/XWzG/yYyv7
G1hL0d58QTbdQI+Penft4ZtgFa4usaXaBG1kwV2Y2NPhIWpG213kETuCYqqdblg7
LBLvWoKXle6tMDeRSD8mQurJfDeJwM9eQFCPJlv06hOvBrxwBiir2ZVuj6b4z2po
U0sM1E15Ril/cFZJbai2BctT2Vpl6L6IQjYHRUPKACmfQpW9aNqiCoD9YVfdIVAs
kGxr6YPE6z2D5/3RxLgwPagUOyXpwcqeyMTSI2qn3Mhopp6eooDVjs0KzWZACH0Q
N1EcxPgRvrSaWngpgdBAOBmUr2Hm6fVQawDTaiP9xG4Rv6LkiEvtcgFQiOt4oCPI
Mx64Ff30htR4HkNLrr+LD0JJJjm62v6WVPShr4grJNi/Jc9f6Rl/nVixmTMKwGTK
dnrjypws9qaF4S4hPN7JNVlPukLeSoeZbPqZdlOILyhHaXmY9tgHGNK+XErP3+rr
0Po5P+5gIm4xs5ruhxMxWrtgynsMGpwOuzigWuGZ8vcLP5x7v9lm2yKZZm1x7bLe
60NExkJoBvv/c8wqlnyIudXB2FYXR8Ub6DWpxMWIlHt+VL0DScb2/JV5HtJdICTU
oAZ+/gH6gYq1qgSL4tKdacWiyHWOVaBcccuUVR2uVbTnEQIbhUjF9hRKcxO/X1LS
ZaPFTu9Y6Qx7oqMmetHH4qg7DRvZljjDfsRlJgEC+UEy7nIuBhZ9z4l5rb0puvvV
ozbyOka9bJWF1Vi7nkMqff0jHjlEhvbTi8ESZ7IRQMN+eGb0MoD8ycOY4yMfnQM/
Uu5YCb+csiIUxIujBLasO4InRcIBdV05kKKO6+miFzbI2xjaUwR3amQHJEhgvzmo
UKfKPUmTkAFeYmEryB/7Qt9LOW6VwxKmvxH7o+0ipKzy4rouuxXAx/aNhRsfzPf5
hF2+j+MWWky1FvaaxRm79dDy9nZCtCj0pfvxWJFx2KKN9dBX5d7w3guRgYlQtFC1
l/BRR+mdTK6kv/nyLe9Njo5C+rjd91I9HOhPpBo8Lq5OSLuqc5R9LnDPYzJLKxLV
4Lut5/xShj2pg73ND+GdgZ2BpMsVwaVVozXQvDh1areuNFvG+Cb6Ik3MnSVQAIwQ
h/Tpgd6WN/UPEeAAaKybttmmMUHaNOt1GkLvH5ZQMihByYNSvYANiS+FlLZpDQNf
/w185iqYWdFjA/wMTsrixfL2HAxNpIuWzDtHaFiLAhcexixhOe5iNBfJTGDSQwg2
4/cUkSiTw/cyYofeAUu0T23l+JIQVCRuzejgUXmmuD86GXAco4PAkeewCz+FM68a
pPZHKNSaQSS7d4bmrGxPjUdKIrdW6eqppoyvCxQo1zoKTQzD6RdtgIam3nsJuI4t
2QecEYWLdygBLG0olrv26J+nKIdKwtj/xT7UrxISE++nkHlu8cAFBgoXCUkHRBZL
DgfHGO7XmPfSi/PdRuCzKsmDycxJR1Jkr/hmG7tIM8xmhbQeFuV/JVx38gEarKQJ
7jgeA7S0O1aEsYk0nPpr+hmauyKy0THfKGYQEqtN/QsrfNIYJxy1E+kuKa4Edtz9
aOb0rxcaAAqtZ2Y4tmQ8kBY7yjnbWfaxLV0AJPzhsxoQhj+bJiAnk2pVbUugIic/
JDAD0vmxydUQkmdMlmGVxqZ9vvjg9tuDRpMIoHsQEsA2BLg3NQlx67Q87kdFnVPS
Fbp1C6wN528zlRbmi0iph33RK/n6fXgxUFQZPcKGJbI+zMAn+iWTjhm5jhtmJVwM
nksBMaOtNNUOcXeXVsRsY3aQvnoMDy5sGz97PudUxwDe4XhA0x7noDmGMZ2G8C8f
n69W6NEbM8y3wyHNr9+6qFYsIn8y43rA70qjXZfB7gG1WKrwmPKAJS8L58u4vmuL
NtzVjlJNwh/Hsf1+FPvhqxrXm5wyR8qajBDtcUfMCGl9H9+xfFM/8G3xuC62Gr6S
zSzCdbmK1VzatkfaHChnPfPU01EwhbgwDQAJALk5ycCYAP2p03v2uqOp3lfSQW64
C5SpJ+GV7r7yqW/b+z5qJf0dxaYDbcKZV7eHEYv97PVZVjMTQLfdTlWVipQiBmjo
C1A0wtPPkZEYhN24QrlRSn3xyPIyutjV43h0EEswOiGvvqBzCyin24ipCteJK09g
eldIbtUD66yYeZEbU3kCg14Vm4CwtO9xD0JcLLKFhEpDQK5mFsnM0RXcqLy0e90o
7xcP+b+1PccchxLepNtD6VmynisJhyCXYZ5XdobXufxtgJpaqe2LeLGKZswz6eQh
NkmyyasSy/hrF38ZroNHfeRR79kRepAPuBX94ligQVOCatCtnU2cLiZnRBwCBzrH
bMgFMFfEqES09ywhVqaD5WuRSEloT6iAPiFef+D1yW2lle0Kr+jYQP6Z9Qu4Zl4s
FIsWitlzUcWoUji+TufiM760Wq1ranb/PdOeLYbSYFXno+PSUdprYgbBOgDg2a+c
hfTgoUof4vg9/FE7IaYcOUD93V4TDlLiD/cVAqyOBEwAFbzRDXGdiNCrbOWWijiV
rFeO6SbEjQKrLa/GMJjZz0VRlExy92tG7y6v0/2Wph/QrBkv+tfaUZZApMdgXLOH
03cj/J/LEszYd+eNJPmcW65zZBE/vmSjVJ6hKc7ZvBxNDD4VFm4SycJBly+moZY8
1K7N6D0NGi5wmMkFWfXKogVxUzO3iE9nBjJ4XCfwmxQjKvsHiOXKwCRglFXAaWPh
Eqx9Wbf1abJnooLBNB3YjUJGWLy7ssJuRS53OGsZN+smBzbcSrZNVWJu/a/S2aOE
l2u4vTRwxZGxeNEIZKbLqNcgGuUQe3HdrJkzKFpNuj6SC7iBSL5PIaO0o6+hmw4Z
OzcXNL+QnlYOefEoU0IEqIzj4c64Ga5Px9oVV00PbBawscE5g4NlvqFEpecyulJ6
HQ7mPRX7Y/2wmH8vMIxbriDcWHAyAFeg9/jSFwgf5pIGT8Hknq/jwzL1c3OxBI1y
UNewfDq3PhvpNZymi6/X2G6JXe4cs3wiVuj0InnS/zUduUP9x6/wI5EEuFNsgd7T
M1h2PmfeAxumJFBh7REFEp10LOH9U97/yKxnhlGplwaK9Y1CL/596ltL9AumA6+X
2DSh2sR7slatQLqzwFRrOZdTeTUcqJocScetVM1QGMwLRfGtKfy5y6f9WXHJV57O
R9Lal/IY2VNWaK8jQWfZli1Xy0ReoDDznDh0b2sKPF5BuE80pwGvAhs/w6OFJ7v+
WCUc1E4dIqd7oF12c89su7ux65nI5hDAj95RSd2125p4dx4SMJNAW4muv/Hk50j0
CyqDovJLcQKAPSkgrmDBnKGSQ3OoAKbms+/SOn3voB46LxUf32Id8zIepg62krBb
7YUauD7nlU2EVTBZJbjEhqbzvat765e+slhnPTSuKucqKh4w9ZQurWdD/98AbTVC
NvXaxTEtSDHaVCp/z9P0PIcvhz6EWvzozdj+6r7FOUFyjAWE95C8FfPQMJdofo2f
eH2ILylXnzX4I6FRydWqZhDjQWQ28LNj7ZwkRYKvSlveXe5mxIx3sKPjwbAE2tfu
MYwk+FQavdYKRQLScZJDtZkYZDD33CZwloWVXFYX3ljB20ixqCEQ1Sv8MCWdas2u
nTisUDWa1CcCdsOxjAmdo4b/QMu2+2NUJszCIcH39s7GAxQasFbnb6Qxcrj/lMyh
0aKJx5zL+v2C3jRlOzbBH0nTuujE/al13PfdmQs6wKQcabnfqbCR7Mkr32jiOWYW
I39f8cSVr09As23Wr1i1BDa/OoUxjonV7Qo5+VpSxPwAwcZFIPiSI0P/BrNmFYBi
WDln9Iiwdb1tW/XPEpo/1f/E/e+s2WG8xZQPPSTYzb0hkOywXDXkGO1cpvgdnHN5
OvntlGpXMkNS3eIkt1ginbalnrnzMQVIyFZcmrkbWliO9XIJ+8cDDQQ49ntC5w+O
c9O+VLzC+vvgvjJ+7ETZ9lG5ytmq/yaEfBk2VO7dn5yy5SIGqSLA/0Th0cTssClA
EnxXehgzO8Fr8lYfHTPAn5OxmhdfcKDATKN3dlUO+0WznKTNkwO6qoCn080L7gcd
AsmegRZcVF1H6ZcV3gWahmIrkebZb7ijLDOnN5jdHY0EVZGyl7/GHIkwiwwxTzTP
uv3A6yf5vccPvxeiRecMDqVnnP26W8g716hC50R28yEVKw3D7hNYhBr1RPrdFZA4
+prHJxmNYR/6uorFz455WLaMNGbaTnXFQoU4dQ53EemrbvBWdgsJC3RVLjZHynqS
mum/rgSqdj4+4BNZKfP5kb1o/OTyYEgdNKs/zkmyB9ziSE4sf4INikD633JsWLwS
SW/QZaKbY5sqGlD2rcRkEO+dIqs4/M0Z2BqTcfHAC10hF+ldgZTUGtp3UT6FaLEV
w3lRl6yA6phAHcbyBy4qdPptugY4d9vEcUrc64/TGutY1CXO++u7TRDJtv5xGg/F
2qxAQSwkh+jJdFN/ozmqbJ8GIx8Vd1O79Z+wVTI0Ab7uc+EtbLwXMVWuTTObNOSz
U+OSXKwMtU25doGr7OkTW4hROA5ic92Mk+j6qkGP2Q9PPzCJETs3qn51LFPN2Pdj
YwVnD6i1eaeWdtyLtV+BTecZr/2FadpVICrg02chSMIRbcsxIXLOxVPaopz1m8hQ
3IfL23hXEjT1t2NX/jihBqPk8RzYAsR61LRK4tbDbJ2O5XGEq2NxHtqFUaEZ922X
diLk5KAaJVplAAB/H4WVmTxQUNdt2TBQ1EUO1gzsDl5xgVdT4sOPGFb7VHTqf4FO
MtDkjQ3yIgfdWjns/qfBoGNYhmI0VU7ZQW/KwC4N1qqTCsmFoDdNkLB5Lh6yJg88
0tBzkz+dwqyi/16NULxBh2wcFBNcwtPh+QyhIejPAEIHY9+6bF54ZPbLExJ6narh
++JfqRLHZUtjaIZwUB0tca+OMPukD+6YRbgjEENAoJ/7WhLRt6KGrCO3nLSlgxSC
LFRa2KGrsWrN+G0PIhWNv51JImnf4/rZWc0lWOB4FMBwlGEM+Q4d9YC8o8kuFgbM
M59D+eTV4ZgCBMg3aYHq3hFJDpiSPP/5NazxcINGB8xhdsHjWkUGEpns4PK0OEAW
jQojyuMTVpWJER3WogZOWK4JhBR7FvtI9keTNk8Q31bHIhN4p/nLOHb319+/UIcW
ThOHMolvjWQ0I26t6nfxL1nIfOVnhLcvOZ1jubxHc/oMBQB1sISArWoCselwtLvJ
SwzUBAr3bvPWJgMw7wU1CwuiDHg3nigI3rCUBjYoVVbc2qzl9w3ipSY7o+fvALoy
DKDOdvLJRTuRXWJXmMVcAbwz7jVYT3CrWRraB1lrwebXWcAd29n+0kaFKuUocoTr
5oSlGEnrkrlBupOc2XRqmFDWs9c8XpI/H6bBHiSOMO9atmv3CfXt3QdXR45JV+oL
Pqwh7iYWKbWRmOxJlHrJOQoCDkwrpw8o+u8aiWHQVyJY0/Os6AX72vaEJJCRhIhG
JoCoxBammCk4SF8vrLhAwoCtyx0nhM+s2dAI37dH54qIz1PLJuUOJ9uKJIGF9+uP
cnGZ5FrcFAZCOk96GfobFz2/sCxBeX9+qQ9sjWnVurPQ5z9AXKRsdz6egZd/iNRv
JrlMvV/zN4jmSwVkpNvxOY/S8aT5SS5w48rRUVJy0zoEin+JmDbI1uf+qfuERJxR
fAmeUZX0CGvqh8bmUArAihPUNFfPcNYjVHTcEkF8uZB7/DbJvCuUVkQiFa+grnj/
y7OMeQ3JehyY2z1NsoxkcXNe2eBe+qOSdASlp+VK1oVwdCvemNDxutKtKi5Ml/kw
x+04QbPW15uNdLXKuaeNYClyQ9yyd9LdgkRTq3QMHXbui4Af8js9Xf2x/CGerQ1Z
NWU9xAz77+H3SUd4RM37Iq5iL3K+YsC/ljag+Lu1vM2RwuF2RCGwD6nn4+JtQuJO
FsqWhBV/+uQb4nyyZ/MbBd3zRZ6YNzy/HPuvCQl5ywyzWYtaLgDLKZeyGzg7zcAk
eU7a/pE7zF765NieJKJsh8M2IKCwt9q1xAhWmPcR2YNOx/DvQxFcOP7z/tSIOhoH
S+yBF4dWhlGEP1EhO1te2Jcokp0PVNFtZVdUk6DIvTaGGn0/O7yo9la5EOA3e52e
dJptl9MQdSH0P1yWC80lm0FmyQAgwvGZY6cTPWypGccZjzdG0ROV1XJ1O0ceIJhf
+QwkzFWOrtiPdAXqsGdRcOu2zesyDaFG337xMMalt6lFqIHHN3YFS7c1bMCbs5ZW
RsoaroL/4zaVVdNOrJFKRvo30Bbqp1baObZ3JAcIz3WM4xHWfLwvkWtYTujsPSsC
OWg1R6LugI+vRpovn9ME9G84WsxTZV3II41sm4WKVGkAzPE1XBAM3sOBTPzgOfKD
DuIr/BiDpHuL3HMw7tiO9oUwnpzMVtqhE8mukPeKSVek9/NQBVmeiIvdxULPp+o5
R47y9nUi9AjlwuPy8Q14MXNQ8KAccpoNQs68F8JZIlSY/usEsnj2DzqkJVHQjrKB
NR9emiD6Yok4WSZy/eBrWnPkmsamk0ocVquHDDzR/1MiekeI/hdHFVcfuLQMdCsM
1z7DQbH8/+XlZBup2Vr2o6Tz0B9c8qp5C5VNxsxFeiwqPagMTuv8mV3BbhmhjFUw
OuiX+1fL8luzeukMchcfcGm+jeWe2F7Tt2dcujg8ZlVQR2S3j397NWT0zcNtH7RA
P6uIdvKJUlM4jIZ6ESVlu5fW/HYzR5/6ltsVNPYdnLKlaJ6YQOqPRofCFTg2/AWi
KJ/xEj47cEI63mW0FF+xc8dNv/qx2WZOHi8zBGDBczeArQ7dC9l+3S+HECX/DU0Y
mfH7w7SqRI+hI6F5yzZjFeOobRAX7DqS2kgX4Z9DNzwSE5wqQCsA8YY1z2F2Epog
PZonTjHcF94JsQMaYRAz1+f3bgg0PRxUcYhbgZ+6210gECJobdIgcqtXWD+tz98C
7oPTt21lRn+qS7sb3AS+yTUojyNmi1J5Jmu2BKScnvEJHlIsFq8T7HUVLsMgAyB/
dRpPlUbElDVZGZ1POXmti86GbfhGVAMPyY10nBWrr5Gw17gZ348k42pgwtTRKNa1
giYqWgc16xQ9VwG01RKEDI6sBHJI2Exei4OUzNQGuCnEL3QbtFoatLmmonbAl50L
FJNx9Dl2UEiMPbZP1RF7ksS4+EsUWK6LEIB/HYBzn8/Meb7CfefAGfIp4jengvmA
Wuu1fiHiv3q2SgUUnibsUMqyIJO5eHEgKUcDV8dn+W0uYq41J1PaOJS2gXTChP4T
C3wlisF0I1YU7m4QZkGmHtQDAFepNDYo8EYJC21zv+p+yHpWYaIORzn4gQY4Ul2K
fgfSJFgeNPLb43U1ymKhG1XTRVCMfTQ0ixct+JPaDRiUeU3rhF+nPeVrJZv/IXeA
tt5zHdchsMxmkoPpAQLc8nN4LEUCHlT74sTeQ+6zaMawz4pMM9PPrGEHy78StogK
lzzwwavbGjMIPL0oY3lgiXOKLKtglV5Ovotdjs4bn9YU4es/P+dRI7rhCPnkdFBG
HC5KqOroKcgsZilKfpe/bX3k64YPZlT1lHQuMSux6Pak6nW91o6qH52VMTa8ySdl
+Lq6RZrkjJCl4Z5XNxlj30c5tswTIHVQ/Ynadj4OCGIHlb3qjMb9B6pYfdv5vua+
HVVGzGEDRkKil69D9+VFE9hJXBRfNJpjnEP44JdRqc2NKW4NBnusEg9oz1c0egEY
wYwxzrOdMqW4DxnkVA4PRPMHIQSj/31NIJZSsjy6MuNw5kh5ksZz/IpgdAsibDdo
h9Kl+nDCBogLx53eumf0VlTbr5duewNovlYk9qIrqWX2ZekoozHn0jKWNXPmqED4
1mjKKstR/apEKd1EgOaYqhJEqb1HqveyfJzcGfJ7BA6YhNwDdTcPqUbYBot53o+N
mdTLw2zPi0pGH5RJ5L5jIN4tjIya6qOdaq1RcO7AAdjprehOPyhknrUV+oh6qvSZ
hAY04gkafyYfSWtcAjy67fcGwB9VZfQiqliSRE3Gu8jl+aNsGeCX24wdIGg0bwSu
vyxpWOljSUFO1+f0XZg5qGy36W1575znsSqKtlIC1ySHr139CkgMT/4RsZmZ0PLZ
LH2LoMQmHZJk4owdnMm/BJQZfwsJjdVMuAH0pQKurQoZH7TDH7vaqPzBRAQtce/T
UuFvJtoSMl8F2UVXX2bFFwZJDTR8AT20fSdsC5DaBokE0loB/kEw/gkOSAgJTLpb
sD1hk2DcBMwrhbX6mJt3Rybf8Ae+jNOLC3LOTJ6D2qDeotJVbEVBhzI12Ip6j/LC
yZ1CxrIsUX7nAJJAyFakdHycK4QHMEKrbfxtvDYrHTkH4hYxWUqxp0Qm1BP50wxu
VGdDtGKBPb1zxFf6vEHND2Rfzd6R2BJ668Iyr36gPcZe06zUgDlB5+7UVKfKj8xg
ZUcs28lnPDlb8Qcqem4pCgSNPabFDtp9ggcx0jQxHBjCuei4q1e1l/84QPzNwBAP
UuOwI4/sNNwUjZBAja2COPXJYdulV5VkaWaWavDQbfSmTIokJoCwn2Tp69e/yPpe
YP3LB4tHw3+/GuzixvdS56fgL0thHKe+61EyLRai8KnUu1rv6B01fSmOgXWf6Hit
mI2+Mx+OsG4JcDDI5vuGQmEV56WU/Pivczb/viffBgP63laBSKjvGS8b4A7bkrHq
MkaZYfg7xU7w49w44TIxbs+Lj1cxWhBi0lGpgf51ybB0ADA6TnZ821TTLNh+u2ho
2ebKzlC58Ym1FDZ0xb1PWLCk2zzjQeBOwdbsLSJJsaamy8KdkWpFT6+jrzLuggV/
OkblLFiopbzjxBgDAFAQTiIb+MEQA3LqK9nbb21UBLWhvVV3aRjEfLVkse0Nas6o
R6Pe52iGL3rFNgR3xC4/fMSuRDEWwltjzPwXvB5lhH1vcnC+G6lT6qXmhXO55h0M
ceGMHBbCE8HlfpnU1qKsLeOHMg3hn53VVKS8LllHFDgARaZgOztOmW0bCT0A6s8d
qB2XVPtjP2LELot77aijrQC6B48m9jyIHErPjPO+w+4e2ZJ/Y9swf7Uzadv4KcFu
XaWlFTnreQUf0c5LLn+mSMZ1RaaIAU234fEVC7VQMN48hcGIHrZKFh9dd6C1pKi6
bJ04Yp0wIQcFp2kvJ6aFB9hN/l5KfTEt5T+iNrRXJT0IjOczVynWVcWUfXIsW8WL
Aa4M8rgxGhPjvL+Hnzjoj2y34fcta4HfFjVhTEzjHTile1EDQvuRdYaA8HOzCORQ
UMkrzpfE6pixnqLhDBooyy9DA38+upFOv0u40d3FbtkO4+JXT97u2fgbDysJnu2f
v0xip3/bwbkJnXSippO00hZx9pcDjuE/Uydn8Zu2XpXk65edikHSLfGc+hv5Cnm+
euDBOK9wl/628kAVbvfWb9X9+i8HNTyXWY7SKVKa9Mw6XLBfQRiJfOQBI/4esQ8F
8ZzH1lK4pN7VWBq8i21TuRAq9sWPmmPgwwDTgKCjtLn7Z3YV04tXxLuq48Dx9ASk
iaagTNxwTDpJVegvYYI98kZwxbj+pYxt/uK0/AUShRkTuFGBlifg9rbWTZD8dASd
+aW8tnFVSX2Ntpmd8fpDboC2zP3kiVrv2dKqplCfHIP7vCA19Dbe5x0UMn0nTIxB
Lvza3cbFj4NmVpStPCPUAqNYgN+Gp1DloqXTH6VZhh2RugGOTXx66BXJgAinrgqS
eUI9966S79rb/jm/kw+pCCuYG9+S33o3Rmr/4bxjCogxfOJrD7clS0djrIT3XwXl
Pw2mlqNR0LPqGPnseL/SPX0DtbEd8bRt+dz180flmCS5bT+BxMBfRhjxuQjMLVcf
GSY+Hlza23ggxd+z8uSQgzzgQtHf8e4AGqoRcA5DclvDYZFZWLPeqqd/ieSoWTn2
69FKwca6ZkBJBGQ3vgJhcoCOS+AVy6CI+y2FYIS+UEcEV1g4lVhTkzMlgJaxxIiW
nAgYo540DtVAXqXM4JM8En2IygSyEZPvJ03S+38beIZL+/gzvlDcL0n9Q3T1XTos
Hj9PG4tMm8BHtWoIqHb1GUxuJdY/7morUyyPEJwB10YZ7ddSCedC05d6Dd3wBIX5
BM/5b/0H/FqnngFMyRLq1ujz5pzomdeEG2qqG+uN8hfuyxuJcCx1nmSFl4jdsCPP
Jq4PqAinn6igZZXuEV3W5jKk0tiDUCH6HY32PAHhw4qFBsbAtsBKtmIY46KDqM6O
EEJrdCl09ubqFnHR1I7DlBuIZUXAAXTDn5ztBMERal//Uyr3n65CpTlk8ShoRZXN
77NKJ1sZ4jo7/BC4Clg7gdIbdDuKA+NKEkDA8DbWiSHp+OTg7Tzp2ea3tbCUauXL
Y3BmcQUVWRf5sKyeMLzIvfApDG0SkUi/PIwOKtSDDxFI6hXiUMK2qd0ZW0F0RNGW
M2GVW2FTfHka1tE5Oj86RjBvUcPwMUWuMNITkFFjxGCNBSLh1SDGX7ExwOEyi1Gy
mBBz9oK5pN8YOwSRWCSJxJT8DSpug0V+hR8+zjI4qLlh3cmEX7SAZ/G8LOlY3Q+8
S0ku+v51nN7mBo0gCXlGVqh1ZEJmKjF+SOU9yJLx3hyPmRQgYugbyZDOv3fhBwGy
TXjgGRY9Ni1uKcOsfMtDjxduuOGLZ495EBdCR3p1aayN1iJMbz78Gl62yvFGSIVZ
ffe//ztAnbrQLGuEgPgFP6UlnPpLC+IEQlyvhy/BG3QniPE/V5ixvSaAvc7FsAYf
XHZyjZx/BKriwi9sElVMxEZOSBRxHAUPWImQtP+n8nC7dKMWfL8i13Rh9fWPuugT
gxRxyeHAfbZrXVY4egEzuJgXJuyNzx1+IrnNro7iT+QQYqSU2DNug91NG2+ydRzj
buQuzHePkRKL3KBsT/0ylQoPVqboU+IRcRViIVIUipO9KjfFEvjgJb1rxMb6aPTs
P7kIw3KJbsyn3QBDZNW+YEhYx4x1FW2otpQRbZXRcoIQ2S/G1OsWzJ9gm3UV3YgB
mfdtzqE9IaeQz8jzV7cWyqNU8Ak8MKUSFUTk5mu4EZAzDjcH5/45h/bHEgnEeyWd
n/Rn45MmcJV7jXvKgnJkDRCkIIqIRjnXLFB9Lb92or5/mGku9mPNeG016KPC0bRW
JXYXsWMo8ZbCsz0eLiH6Hv3WeU7BChdpG6ek+Sc2WG0OPKgjiJeFrfM8A1f4aiUH
jT3hcZw17e9qW/ekymmPrkhaTDrIDjec0xjJPg3MHOC76i+A/7dzChKmj/jdofHw
sbfxot+GBTkXyBgBpqjJUMAnOX1bHT6A6gi+ehd1op67saTMX8iNuKtPlpPcKDuf
VKp7gQOSV91WrIUnP0gDd9rTHfCBuTQ64tlvSP04wck8yp77Hx1w94vym+m3XzOX
Xg7u9uuixY61Zs1QQJ3+Abhi40cwB8Y0kIAiL2glojVS/cdhBIGQBEHFaRtMNCoF
aCSYdG91BE5hBx2OeKqoedkJuuEJZKafHF8Q05s99uRXWAFUh1TFvMplWX5uetz9
M08JieVvlaD35ldjjquzDen8CZ+GfecYB6AvHSm5uZ6yd/869ivCxvx1KhWHb3AG
q5AuyqSIxNAg6hJTnGPIYDJuMMiJjkHKA/kdPPHu38RB5kH/0b99pUXlu+eBwC89
VXikqUOitU7Quo6b4OMLDfswfvG8MA9rNzBnAJvx9JTDWpofztN0LSftFeOXDhnq
cyeb1Yhol6vB0mVasqJllQOWjixkJ26srF0PsImQym4nULHY0T2Aquyizs5zgbIi
3gX8hrlR6iouWxOkJjIL015qJuc54qQa54xIH2oEImar13uIrsjTKxmgsH5KEASY
JxEZfuLsdqv77SaDP8wiygVp8vflaAtlBGP6jY/caJLriAYskib3Yp5m8SSmQL4U
fnGF0iRQYzfZqCsFQFWo19YSktxh6+/IPZjBfJywxmi0QXdbTyV1/iHhrWRCvFJ8
w/5R/JVuyLUzVqc/MI33hyZPiHBGTSqIofZQEp5aaM9IC+s3PWtPw8J+sDcTKfB6
BaDLKtxI5TetsDcjJ4maUmGEKLjDqlFjLptJraRq5vreGkyMksUMMqsbYMB8J3/F
7StxIrENwBGN5pskz6RPCPJCVLRZTNB3PlYTj2MKs30P8lbCKO/ViHLQW6C5Ywnq
J6BYdTfQQ+SSrekVh1h/EjhIjvNiqjDqJlj/uL4qce00DB68OmACWEVpOZRxgBvE
8tur1vxD1cvhaOSELRh3n6I8TMzxa62xhHwSWJEek3XVSRuom2JzlvQDKUyZb16n
GyWcjVAdWIjwsbtPS69q2lt9WmoBEVbE5NqRoXOe90zyx3f3Rt1gfeIohGAlrIF7
nMU+8fzLs2ylnN9SgvI2Otkr3hyXco4AifToFxLPvN8bev1DZk7ahvRjAHNgY0z7
L6dRcxh3Jj9ye2GFa8sQ13st5jfbhtUbg0M3sXQUNviXCKPMwPr+o6BY1xbJKSCR
MJz4WQYZoEX7KIxysJHB8I4Beyh1TgNJZLJDpaDze1y4LEpVyNOEHew2IIslzk53
H4yXPR3nOMkMyg+3tJdtgfWW9vRjdMFlGmMmgfSVGmDnxUOE4hePwktiIf04xTww
704WBLCuBpYbDr6NduR3bsjTIRd60PQkdTrAysvv1LZ9JsDQSToVKAbQVOy+gJJz
owMlfw5BLT9+aNkPbMdrbBLVBJvjlVrCifi/bvS88+lXZe6hPVm/ImwECvbISqdL
ILVy/O2wwOxrQbsbdHwT1z99ARYmwg846JLHfq6yn1W0W8zU+WJhMoglm/TvBZlJ
N2UqdnVN8B/jkg2CKaPV08DYsM1GCeIK2/bsPzUb7WXfy7Nbxa4f9X8sw5YJlB8V
IYv8XRbrpYb7PwXvQ9YmFhYcGgzFzY8uJA8x9NTKNVJHUxnhBZv4aUyUkH4uSoyu
xxKQUBa87kxBWUTxiQObHw/g+44MkqqlQ5vB5GRkxdfQSva/ZFkKz9H19Gb8VkY3
tGY7eAVUxzpNEDqYctIvAJtJvf62brESuNqRA9AANGRKI102A+R96C+0Cv2Q0tJh
BQQ7FegImWOunU/q00PUfB73LhoaiSOndv8NWhnZHtAaetsb65muqxra1+WXm2dO
5A5tm8JoGDz0IlnAfARo3QG/RJLuf8esvsmpMhfg7MIj1QeNZyAIljJ7RslsEVcB
BT8/J1jOs4fdGtzYTkqLEYTi4VTjlpP2jr9yqab4FYpP3yMgKac8wdGJp3JGXsUL
uYZmv67+gc3KbvBK0TFRMLFKGVKhD/IPawb1ZjRjkWrGDE643uJTg5JKqN1nNdN3
7f0a31cPFJOztJdeo3R6pRQ1bZEdTxIeOfsvjS4bjK2m7kxvEAZ6OXn2O57yi8TZ
LT9h0+ScXy9XfXXtr1f0UH5dpAXxno3C9FzP93GJSyMQP1rlZCJgNccJqAZ/8E08
LQFF0wTIYQb7aZYBo3RmHp810OXK7PwCmTUXzd9w/CET/9nhxELvYHMA5qWJ2c+n
VXHExcqHNmH71DjYSt+xDELvarDcGITkTHcZCySPa0PpVqFhXXfJRjufBPSTvx/c
tgDYnnJO+HKvQvx4n7loXqyZsZVscRNwSzSXDFrEkitu+5aJSnhE5w7W6jNUiQNL
t5oTfWwBDfJM3JNoLdG2Qnm5tQSxLHZ4VdKEMuhXlfgtRKGJeD7/qhhw/Gl3nX/o
KJqb7ov1JDbmGGNXkp5FtWZ6MwTgXBXPkX7kbbAP4gJQ1s1gJUWlD/WBj3105eBv
kANzMedHuxbL9rt0+iK7gvn5GfuHnZMshmfnNQHsrr6bsEdVaoNwoY0jgRNzAw5z
h6fPgr6n53dsKTQQgz9bbqmKBfJU+SjMW23yfTETz+T1I+161CfMvFVinAOWMOC/
YaEDXO7DHFiTplyRYkVG+vETLYk2p5jZ8svQLcf67iQqYxLkKW16CwhZr2U3cE3a
mVBa/5xHzRtiXlwsbZWKHMwqw2JJ56Oap3EMkT1Xk6JD196b1JTdLOQj85gjE63B
BHFfjDSHtTH+srO6j7TKsbXBkyCSg1BYxH5HWl5tQYnx+RRP9ZAmCb/Ix8QGLyoH
EgRlaB60p2hAL8/zh5u89Wfa1Ti8VTuZ5U4PBM/1TR2xFFOhLLvDF4O4MTa1Iw1m
gXa48iWjklVLySnOjDJ7ZMlfuw+wdWgdhL2BKTQRyePabVAIA8Q2xcFru/VxcPGy
AYWzKPmtEfR5T4EPrSr+s+wJ/2WkSAWlZpyWcUv1VSUxI55LExYt1uI/xKyu+nXZ
yqXGu1yOk98o2ggQ5frjVeiIva621+lwpA4aa/fyuqtKuiaPEjLgmo4h2ucPZBR9
6bboU8NMikb6dx/jFwmBMJSJidZs/2ELXMPT+5CJLovn3vHFH6znn9IZDddGi4Fh
VnxZnhWK3VyuoL9wRHDPnlKca+uX96Mlw2m6b8MhognLeYGk0UUy/Rk70bFnLrqM
5sT/OtdQOoyaPiVqgmJGNSJmC+loGYW8pNheWLtP4yiAXQbIVw3fujmPMlrHuZuM
wqGrSpLRpIAGaHMSkLWsgtWAhUZRDc6kFfZ3vLsQXmjRDPzVibNCFDR8qEFJKdKr
KSr7hQbCny7F3gYpyQkDnzLndkVHn7acUNeqFenRwONraYQgDPUBNca634FnQHRf
xUUXq7uhyTzlgdgXNwp+dx+hD17knHO7j4RXZZmUre9OkpWHBCWbwWVN4h4p2Dp+
3tuwp5jQpt8RHol20Ce4lpUDNJqwZg36XqhlA1e7FhNYzGSJHTrl+SghBMG1gLqR
sEvqXTsxWht9mhsNBE/mrFysFSS9ojfzmsIUbxWIqXEXnPMCLl54xW9yeE3W57s/
qmPm5aRnT60wPkMK4XdleVgXJB7YtGXWYjGNRUs8kdkRjMn0SPcFO6icSZthhcjr
scg2FPl4gQHhzOOak9W8j5Qcgc4CJ+EIntqW5cVM3PVYcEuSvVDMsAMcH5AW0uum
/EP1/T23lzklBU7fQF4cM9e8++/Uf5v9lgxW8NKsujPQhsAaJn5+9zXUF7oca0aj
YhGn+uBDXPHvRacs6gnFWy63V2GgZAHX+NbhxCKfERaCm6S2pVSMaj4rtfeDVm1w
oiWdah2a7ShkdoIKEYfwGIl/AD5Zxqj8kzuFuaU8jzC1bEUSu8dvQD12H7DKtm3v
3iwWz4pECLkUmfvf181G3h0ooKAPbsLvPBhsbI8CgB7ylpAkyN7yq0ZeGiNdCG+7
K654c1uhtYVLrSgc/EDyvDKGaWk1L3oV5tZyOn19+wqP5A9YfmdF7jjxZ14v0tI8
GZNokHTg921Qm/Lwpc11mSPCL5MmWYOeIndLaHh0p8kys18HCU2TGJGEUpkANb65
TjspCxVBfyvOJDLpvyWP3ApmZAK76BF1Gn9Gyw0z7nG5Wjr1sfwxuYPeHTbXqS+U
QGTv2bUczSB2mI8+dUJxlaU16GQ7Xj7EShQl9PriyojSKKvDVIWaqGnbaTSwb0MA
TPdFnLJcSrC7yWdTuHv7XanG0LCwJUfJTTymrbASGhS937WjUjvLKMsjdGtVrplC
Qz0f67vk+c6vKGouFAQez8TvIjtF6Jz3OUf8wYGRwr1aoBE39VPAiVi9O3+pIERI
Gameh7etEfn3qlDq7+gCMoQMfGomc5D+1d1wJw6D8mxn1InkSnhMRqKyWWK2P5zE
dEPLgaaXvxHyAmAsyDidZsRooDwMx66RVIWbj9RkpfpAkxHVu0M0NjpI+pz3DSdn
v5splqH8qAi7md92ICnCtGAxVZkg9fmUvWOVnO9DwQt97dYttdYNcGUDQwEs7K0u
V2yPtu7rDqKA7W01X7HmJPSIP78/lnyoNxcD+mfpuDH2j3OGOY1AEUyV2J5WQGfD
udITVbSXfKgittg6KUCnnbnGKtA3wCTxRyWNPzmdxS6PPO+VnbM3WJ3XaCdt+dj3
bzVm/yh2bX5m5djvpPn+kxAHoc3FjIPhFvzlmkDMtYd0EzjdiuxTir15Q7SlCEBU
e4sKSDmTeYNTG1meDJ+R2Xu4LislDrGaXZtKLkO8vMlvo/Be14Uyu/T8SgkPpuTT
YCpK/rDu/JJvw9lqkDiY0uKlQfBKEVNMPmeR715rz5b0hRKAbBZSUHYBqfP3Sybc
/oIiGVjTf0JG6qutWINphcvcFjCZfwI8lGgNug6yXeKnNLWXhgrdXyp1HAci8j65
zzqz67eitZ8kIrqjQMbp6kTITRFzSwtHtujnr9LpQwqpJ9U7F7vF4Xy5hzJE5V7k
bNVHFWKo+BMvMUovoKCTi8UmA7m2y3+G4wkp7gdwSLqMVTh/KuejWzscZRbtHK+g
dZESreL3q4Z16KG3q4nn7DPB8G2iLkXEwakETw3kaHMWuxhCJ2fvD7isDg/WXI2G
HScAFA9r59BEcfGvsfH2HkwtC5XXA4FGy3fQmFxbBH4X4+rD8l3ZkSJMkN7V2DrQ
CyOe0NxeX2QG430CRLfvooOe8Xa7i07FZJUIxhHcslGwGBnXTCGhTlQZzD1py53J
h8uCx8P8bDl2bWr0Ipqg10dI8iRPy1lepChZXHEPEYiDqcPOu4t8DoDUlCsjhGQv
lidgEhv01Vk0k9q18yAtvrf+Jkm1BMw3TMqyVJqtmriQfsufuWzNJyOxj65EC+lg
P9NmAL0pt/5P+lbBJ97pTHJmcI6wwbfTbfkBV3AXxcEj4PdeHKMWmo7jhK0PB2eU
+f4OT0oqmYsftav6Hm8eEPWoUyWmWowyWgvZ8cKHeYB2IlHnThFhN+73kjDzEv4V
hWiZY9QGaI2fBP0R369LzqlDErmn2ZXnkbwEtquJtAThdlz+vp39PXYeYpXavefM
Qg0bb8Bg4kQsVD3DjEHfOq3ueXbDEa1G9wGugY4dOXtPj+MYqKPRa3ap0tLwxQ3G
WSXmVU9ZlkD/OWQTjZkbhZDEFsf24LOfngM+xquR3kLuShESyjeG0uPd2ZaEZZT4
XS+wjH5TJ7IlW+vKqtqwI8D8x8gfY0UqaDbRExGBDRBIC1v1lSbGqiwwHyiVd+qB
5WfUwSAcqZ9QHYy3rpsMhHmxBB3us/QuSlnWXgRPmEwwiQd2XH44uTLap7hqkdJZ
gcEXo2P+F5h5XiCERh1kBWjb4joYxEKO7Wal7acThOBcJTNRv+IF5D3Nq3HWApJV
le1IxiNb8sjhmN1M7U7TRxNQ1Hx8+WhPScL8OP0G1EsxcoaG0wa5slOH/oSJ513k
x8g28GZnUFp6KdCqU8u3iaLzhM8VIUyt1STgifCViu9K/X2oj6WHmnutcxSO01p8
4ZnLeUDAdweHAFCerDIVRI/Uvl5s1y9rKlWF8c6Nuif0lBaa7JiIMC8z6lBh/431
/fWXzp+Z6Q3pa80wmmE35P2TT+VCl8atRIWxaiYEU/ICFYxY8ZBEZclk8YyLy3jn
pGZyXK/RiwJvGGzmeuu3DsyRNPMv0o39P+jjw9awe7n20X4w4RF2p7L2bNvpyXJZ
6hv19RCFgL1gVBT8U84imFOXD0m2T8RJSg3VfmsSO/KcamuZaH3neHTGzdGn71fs
U/fLmkaMi1hpC8fHKjevYnoe5FFzCK1FkC75Jc5bCmDz68yGpWoS7nSrVsM3+RoK
4Jbt32LNvDStKTiGszEX7pS04NBhLb9JvTJIx1zeRkdY3YxcZh3DiO/1xnQa9ii1
M58ck2albKDV96qvQY1ZKeHNif4L6/sqOp2D51oE1PaHQ5dJqEJWeT+ZG0QtKJeM
bMCVJclY4W4X4xa6LtdShiBe/kxQQjMQ6h1GiOeuiBecVrzqj5RGW5mnoZzUZMP/
r9rVhbRkQHhHqNBhTROazigXU1Jp68AixVo8jjENaVSSARXEMwEd3faw/f4Gqvst
Afn6CI/3stp8IeayApJKAiwDlA589qzKWjZUDQPVgNwYuDaeAGgbbhk2EohLUit0
pCdUrQQJNPiZi9+knGZH84ov0aYLMb2gb6fksfpqDgakDDp6O2ZMAB8645CzBMsK
Djx5JjXgO41IL/5t4+fBfhnul20Vhk6xv7DyMzp7IsLoXhQCoPYytYjm11QlD0h2
jefcGMGl3YgkIee06ULbumYIdejHpjkAdtBp+qkbX3Tz/tINkAashjb9D0gxTrA9
ObigUvHk6h9fPUKWNCT9TG/hQnK+ZZrnG0ghBcq3oBPu3VTXZDWJt+ddsL5/eTYJ
LeVGp0KW5OiTAUZkY3EhyEmpDTsCqrJDjD5CyuQZMZmtnvkaQlc+nzga2lBTRw4e
8n3WPfEycidw9NPI9PBjRXfa2cUKvDXD1e76Iv0A4z3gxbE3nbhsNT/HgKo+A3Rd
GqCXpMZj9gnrt6X4gfU66F+9KP8Is6QZFjvUV66QSsmsLYvhCQ5Ds+cCP1TU6uMQ
hyJISEgjx4hHTMKRPsoIXlarCocaBT32NwyD6vXbcBacc8l1iNmGTFzbe2TsiW9R
i9XAPByJ6jgUbSaNkCGHh+vWYt+akEIXEGGngrTWMqZKACrjDjhYi7BFpwC+zbor
Kyq6l9jjzPAnT4Q7XI9I/fUr2Rp+PHEr5aZLzpj2NT7BEHnS1u7pVkqCCaAIHk80
JzpxCzseoAxPoCn/lnE9jfpO4hOW4/2fPbembHuEiwueO6ltI9Ixuz8z4gP4F+GP
tHdrIZBmaW2luA/pL+ZKHXPxhuNGTcjBnR3/cboCgU8EwVt9nnsE/EEVOYp9lzI1
podHRy9ZyTay9OHL9G9VJYozW14MRNRngwAhC6pvBpAtoh09cLoKLmOMmTCd/GQp
hFqtQhNaKXmMQroPgDk8/LAGG/tLoSL9tBnc70MwAnrxZnot6vr38bNByfgWARf3
jQgpHKHmWCEirjXsfPWUlGZWmLS17c9KFNFf4kftd5DS5Jodamtds0qsBotRTYJ8
S2+naZ1yssyjIoNBR9SlxcSqke0FctFACsnRhtlhmKnsyFQ1pyJcks3MNwFT8SKd
ytulOtmcKfso9YCjsjZGLyARfK3oO9EC6ZclTVmtAdckj2gXaj5JoQj6dzmbJy97
cw43X9ePRtVw84r9RU+dTx6UfbW/9KptmSOq8cE3jpqq7DP29/+SlDeqlMeM0skR
dvJscP+yeE03cOzucidiuoxlmZQqzvQGSa5EvpvuugYtixbICELzBB4ktYo2BOpP
n8i8wTWi4AK9504KMyH5FCc8rBALSU8daITg8m4f/hUVRpdF9+kGijvG9ANZT4V3
U/c3A43rfhqee8bQzQA+LO20ao324lJ+wmfxnjV38Wo0QmEMWmivNuFcswnPYukw
zbbPADlvjgyh4f/ieiVmlFo0lawIjORBBTEXqRzl41RQn8Xus1Q6PfMPtfa+A4Er
lI9nJiESAJifq0SH+89pDVtjc3wrxAnK0zTz0rZSsq25zP5omkVVpm+KNsKgYKqv
SztB2kZ5OwE7REIaOIx2tklZSnhiyyLuIgWjoLUMBLaunRKOsSCI8JDGoKGJWzAO
zsjI0zWXW7cfOJ/aVMfGBPxKzKeMul2HiYgDSk8K6Tom325XR1fentCeONyaFT/B
qDkc1bxhYqYFap55ZAG4qQt+fkOh1M4pHFIM/2pVP0pmrJQ1ONjfOiiDeDN794eS
xjZyinJMoEjGW37OrHHNr+67Y3LcARq5tfX5mhmFmXYCF/YESXDA5DHYhOxM7qNe
LwIy8jJKUumS1AozjY01HVByoFqXXY27oDg3VVBOqesLrZKs7nhtVC2pmr01lUgm
HhLIGzD26ceAsZrO5mOEgdCZ6eZqiFPC2MSyK5jdRnCUPldxPDgWGidp4aL2VbS1
9FOjhFgBSpI6T+9o2p2UrlBNMJEWB1pu0UGjOW1vZlQvZak2OaD8MAPVZgENmbr2
YtueEJ10Iovb0jPUfeIA44TqUGXEiCz7uGqavemaLnJKKUKozJdzpB4FukngWGxh
hzk9EX5a+Cm53Hhv1fxWw5Pp4wR5uydDL6bqvIioObZWvFP+evvjBVG3R9Y+Jnuh
BXD8LnD5e4LawWKQfuaqhzlpY27NZ3NAdAvdQs6/y6py9sjikxA7iJyoLvmsA4zt
sC2OhjThwcZ71GcwSJGq36PXQt1kYv+olvP+z4YJG1D2MVTPz8gvtnJlBpuzOKia
c4q5/niW3GxcwL4MLeab7oQNbcbpZqW5vo3LMXNrHk2iVDauxXyjM2fRSwbgkLtB
7+84Qq/Z0OsLdAE6TVhg6Um3PG+645te8KGtYGB6CVwR5Z9+apzQXDBNl5cnseLU
LF5eGM2EAclR5EJ6OIXhdqHu95+4cTCx8MzPHKrp2JvZBQL3LNNKZ1m3EgWmQxUt
PpuAT2m65hu1GrW56KYZGym1Z2VK9M29YeViOCzDChih3XMT59b26tT4hS4wUnPC
cye2YKa/VAEqxeoeO0xw8s7FYjxCiiE/5MR9X/co33YmoRDPI+ukQoCRE0Ynr6wi
j3nagSjIQI7iK5H1HXfChTwADBK9lkzrHU6NmPbdx76lg6s0bLv7ogG9vKX0hfdq
oYUcFhR5g62VzvCd+mf7MoVHYZdS3S6RBwf7YAGgiiuEvVgmq1TJqSClckGLhoEl
MF/3/vTWq/CZ3YefKN4pty0mQcxlRkbJOtuoLNiFquRXl2Y8qVPSurpWXFpQ7GG+
n+UC7L8eeqG1ObK/bEcsaR95XVDFmFXbN18rdBrkwxWv9wVpzXWsrh0RE2bXr+Y4
J1FuxNQP2dFpIzhHN4N7/pFM0a6BbcMVXf187/gvb+ih9oXumG1QCIa4qNcJTqyi
KrjLF1K16fqTMpUueD5iUZCF0Us5IDn4z5/wywpciZA83Ldvm8yiI7Boj0ptdP4u
VSCVUVXnym1Q2J49k/aK9Q5fxz6WFRTBNIMapjkAgF0cYC21eCJG6mKMEMPUesY/
P1UqZUdpcc9QWh0qMQsmjD5jdNIn7gPD+sFRcWH9zyoj10Bcxq3NlE3Ly5b7uWCs
i5s0BVQeG/kMis08X060ybkdOV23661AMvpWvibK9KG4dTYqfsUZckMiyKHhPDCh
abHeRGlFs1QKxzG2e6zcEgv6VptDE65Uy6SIagmDNK7ujUcnYmHfn4DklXuLsGB+
ZMsWEC/fDlhzp5fb8NrclOXVewA2WzrmXHKGumnCGqQ0I4nDEG5ThTQ6e4U/GLtT
PDSZTo4bgeCcOW5MPzGr5FocUQOOa4iPyu2vXplZISOZdy51Nd+tC1erkc6QbLzT
Qzv43aVVXW5HNBzarjh6ws2Lxe8jGFec8rukSEctKT2fHpOk8TRg2kTTH+emSKal
ZL9rfvWQf7dPM+mDc38P7xdLRLB6pxcZktHTOq8NXhJ8/kzQpbc/nvuNc4lWAh85
asms37CazLUhkOGVePY5R80foR2/cPLCYY0HZM4+vlr1iQwwuWMSkxrHATRxkxpV
XWwSwuoxLFufQxN1QZYbSWGqXGookpMI0jLv0OdkQRxqPpQcvNzdOdatB1GXcoc7
nm8Gdh5AZ91gBa5n9+Du14h5mw9SS5pCaPN3TkGxnQXjhJMrE11kxLCcFzp7X01z
XEf61soi9KjNfvgRfYhGSKi/AmpXaSudhX385bhZKD69KkkZNLpBM+8HFUtfxmLs
vjTJs1PoTUkrtozbAg+g+2tz5K4Ye0SAtfNO3OScFjfhNimG0SrNnggM7E5rKW8q
wVogQLRt85OoSoOZcKwqaIoAGdyZxLC21xMnu6Vw4l7NZqcdK4dyBBWZPFcrjEZW
vCbnZxtJLJ4Yb/pbh6XU9feZFOGdbqDy2q4Gf4GMgFPpKvHIX0xeWmijA+5rNrJe
2algA8Yoh9Hx8l8nNCVHGFd8hjvBvZ0Db71gpGCeWOu+clARuTAFIQ5PbQLE94Iz
acyhS4BLnqTUPaEo5xoS4KUluhjCLseh0P9/jgW43u9xCrXypwcmTM2nYFY0VZu6
Oc1r1Soa3nRFrtSvCSeQKLXrfx5gkPxz/9ZrrZrSfYSVOP5tTdiu+HZLjNkpFiJD
MuVNoSfioXsQPQ4DuhtdxdkPVZMhZjUjCvVxfXbtUpC4nirpP9xX5lijJGN2pT4v
q2xGoCuR4C23WkeeofaYmOL7Bu0Te21aDCvY/Oh6CZjS7CVEIyJ3tDrQbqqi/QpJ
kXNGUGJod0Jn2X39mkp4DrqQOhCX4CrgrnNFvo3SXWTQYT1J1Tahu3b3hZdH0PTp
wS8zMlhQNV4magvdXvo8mMjweeLjzPYipCBLGak0MbgcyyqYdDNYfbWOiiBD/rfw
0wGve67G+R53jjZ9o3POrOAf1n92XxLg3gapxv19af83fTIkJarmy2cagwV3LWBK
GN8EaU/UkoCuBLn0SshmkOS1h6GqV0yK7BvZ862NYp4a/GMOX+hh2m0hUVRtW6hh
UiIsiMaoxEAC/voH3dLAa2f41Tjeahj0xUpZx2pIDw9lH7B9OqOil2KiSSKHX+Qs
PH9Y/cMB9b4nB8K+KCOipe8gSyv3foELBz7u+ywSsACNK23PzSxVcIo5uykbrKZk
E26x0gVk4Pj0cYgmOFxzj9UTKeAJxy852cslcavILcFZmOATSKnZ8peMVuOtsDiI
hEBGmUXAh0LavFD0jTPOaxNUk+7/Enj5xqdjTPKyu/+UMvOnUCqhF6udb5uRc7Lz
dUEZk01sBhIQBoJyhO2cs+/DwNoXv3LSdeV7QiDr2dU5/TiVW141sHrCCMFLXU0l
d5AC3HjnPy2d6eAfLm76ERyxlZDFUudnchS5PNb+k0pGH4vaWV2+ra9vTA9xpS0s
V0UEXBO2OkgbZ/Bxi7kk31OGevnq/AZYnnTyPaV7qLB0Eamwte4SV4RgDEiX8FsJ
olmOTOpN9zAgpIAydqWiMz934o0VjP++WmLf4PZs8Gd1bf4Dxs21Zo0BqH+CiA9o
OukceYjbKzuCSe0NQiBMcbpqeExdkc4R81C9EMWLri2UHNc1Lck9o8YK0r69+OPP
+hcey1tOagN6WCmZBUNhCiKVy3xa2l6EHk3poLBmzpfnhBVKr19YDBVTKF0rl5Oz
YBUswvL/ZKjrwlo71C8BIh/lEfAaX9rDhLexwuy1ccQRIo7ObhPtXZY0LfydvaOb
Qk67soJUjUTkqQSbX1Mwe+SVR2YmdlQzzXAp9NmeNPhr2lg5q5q1L1p3xsEG8hwd
CsMJoZeS2srfvJzyRLpkG+WqS6EeVozdAlT88TE7EFefaJubD8d7cpjLe1MFjDKe
zSW5T5tGxPdChpfrBgDz/y+Czmr+G1HQSbujQ/UVrYqKq6Yvu/aH5EYUkMsZyTsD
ygDRtb2oaTmaowLd+bDl/SSif/hCRhamk3T3WZ63mtockq2BzZiFl1+zDcJeG6FS
js/OfEOU3om+JKsX8pzw+mdoUq6yP7ahrIylw7p5BJJbN+IjKbHwMx+XRhOEy00v
lNl4l3D/YGhQE6cafj91rWG/39tezXAYyfWGqo/qJ7JdL9utmpgfG/I84J0E/4CU
h/aPv/Sejffwhm7qKCxrX26P4UB+2HQZBbJ7grmqEsnm0oCZA/41JtcWfAi/qco6
oIDzQB+fBFkFHk4KCEGwuLOYEk9ncevzoNXp6w6mZMz/4law5gGcXJ8i909Gpq62
/MAciNPxcvUEpUOglKhICpC+mySTj+hMsT2OlHNpqBGNrYfP7GQnBbMyrbP7r7KF
EAegBNEckvA7VTU6kXO90CYgmINVki7xmO+TFLpa/MCTxwgrC31ATlZ9R30PazmM
dWuranIO74APeILgRwDlrxMVKhahvWjcxQ3zcoQ++AwcUgq8f7vk3vzU4gdqogHP
0mWLRIKk2dwRUOD2a3a2ZBcs7EEZ0bDVSWZt1k379zzzzMwwxojMuIrddoLjjAth
Zv5oFKS7+l4Kmnj4S8ZY7sLBjGnDyoEmhKmYU7BhYhbgwlI/u4LRf5obWlNn8jEq
jP8e/seVLCdnuVQCk5wjezibYVHf90bgh3ojFaHJkgtNFnmzQBf6CNPkPeuJTqrk
QEsEltqdrCNmvanVP05TAM4AIqgWI2lIxXVATZ7hzO5l7D2CQSAQM651Vp4i7mPJ
N+IrU6MKdaYzvX1b2lm+qOqCa3bW4TRwpmb9SoCZsidQz73s+CTrDgjdbhgDEx/E
qvocRVQig6esK/kTIL267S8qMP1/Q1fbsRnYXiZwKTPW9Sajx/bYFSz2MNDxlyA+
KdZEkqY99jxZoY26rXX/jnoDJ32GjZaRGaVVizhpDjTMha7n3hD2z5uGoEZkXPV2
eLbNoqFEh9flEQ1NMVTi4iw51lkuM2Wk5Wo84ITYRxuThWmjm+GgmWB4oJR905Rl
5MZzEvIXBhSU74848aszdomelVdAFkD5hr6fDLlf1ukM81+SrqilZ9CbO0NjaILp
jqKHTY0ijv6mBH+YaT8BM/Ed5gwZnsKsqjSQDaNMOCeUNoeBxPrF/Efb7PSzOa4M
AHoPFtyRo32eVpgQDsSKq6FEWqqcEL/4+Z+0zrIH5Y0e9pLRZq+tP4531JpBSyGD
SOQ8xBC8/gaQfhBG38ZTIaCO7wulJxJMAQXC9GoRfh3NE8rccgh9dU4eus6zHuXt
NemSCNkjtKrJwnjkFcY7xWwFyMP3GKqK7c+Z7sEna8jDA/zf9MPYdYbunkI2f+uM
egTZyCigwg0miqZ55bWWKw2gep2fA2b6lPRq+arLLavFDOyFYvgsA0ArSxSw1tcI
6erU+BS1CgIYiujFbvsXNNHUkeicjfr/4MHCsJanx0AIyvTY2WRQTUSO2AOydQVd
3ctzMWCCJkDuhN4lSsRq8ejE2et6x+mwndffG0BbTz3TzUMbH1RlfiTiopALcMWN
YgypMOV6DYBmGzZBjgCuypkN3lw8aqD8+lle0FajzPMGfIE9oF7zI+yjV0UlSWgh
rDePTmUAZgySlZlpkLLpJp8dxUB6vrVQ+kNBQC0Yql7NlnJ+ijpaLtb3j2XjKDQ1
ISNf6973C3e4+Tds8x9IvbkHh1DS02+cjZbpU76xGCanrMR2ZQtCLlVhigceipVN
7/rdN/Gs3Z+Xy/b/noqS7PE3VSxBCAs6kG8qj9Z9szjWjnNWd2x5RwsZ6gZgqeRZ
SvtpumH+H8v36G1oSDOX0IJYhJt8XcR+tqM+wlwCa+CdQSxkV7hQSQujupeZARib
O0mWmzrvOIbBchXoZwaPTMCODL7YXKT+4wY7xfpumdLNTqX0jj9uVaeMThqRIcLG
eFj6Lwchiu4hCMscQYANzumLgzR1rtB1owj1NsRYfUUFZHvtrbMDsTzz5umAIlau
7CE5DfYhBJDJHVnQstLfZucwo26W+N/L6d8dSO8CR9Z0A2BJQtBtyP76ItvvT3dr
oNXMb/q1O2hxlEPCc0NiD1fY3eZANpXSefLcAnixDYiNAtRTIk+q8+vDEjPx0nbL
7g2Fgy1bxzwBFLHL/LfD1mvsxedIz1TJi0tCoGThfsiCM8VmSzowmZ3yeXWMC50D
JGkBsxCYwSQEtiTNvrt3OT6d/uDGET8EM8gVoJDFMI+lwj5DDRjEpRZI/JGwamr/
TIosShBDWH3Ee4aqLS5bZbVFhYm9D9K4NajRFY7JrGmb0f64pkrQ3+YkJJBS7eKB
AHVNMz0MKIfiAhqTjbOaYW/JclBNsHFE9bEP1fEjpIcS6D8Y3zjcCKoFsT3OO8VB
li8ron470ZY/qzf5L+CF+kei/K+zm14q8okEAYIm0zFlc+wB2UQjfIaMZz3l+drA
xma0J7XeMAo4AzbHVtf5VGewv0DndA7U54DM9SncgJi6l+gOwqKo8AtWNIZe6TYk
6NfzLFQcyJx+f5oZRxJGyW6HccA4m8jgK0G0zFNbEJzHlQ2Bed/7xxSJcRY009gM
78H+9sseDl9/M9cOlB4IO1nW+GWKgvJpKxRkHzJO7DtZEQtVWTM0hxDja7PN3KKH
4sCpwDzuNcADYAquBicZyMPLC/6yEBLu8y/8SG7GXVdEYr/taYo3CyKD90zxoIoH
P3fTZeBEZDPQMvl9UbIxKj14z5SkNPx+Bmae4xlTsn5Q40wMWtLI9JyXGQQH9ZOU
MgOGeUS7zmToZ+epQEerNmMysCwRvaKZ9u75ROoTNvxoR5kcAfoCNzmXTy6Zi2cx
57oin2OFJUwRDgMzX3XwhQqbTYOjZl0LbUAU4XSmBctlWzIksyQg61zTWorP24mq
+Op8Vfr6oVPmevnmT1oh/z4lB+M5PwdKJ69dGFTMwV/X51y85iSj5DKngJTZa9ZH
Ouqs02f5KxiqIi6OT6OiEjKQnnzQP+hlsRbBiZ8wv+Z2VmxnGOYZJbvNWKshrzFX
xlfDAg3eDazYxICfookoUvdY9QiAg/OLFaxd5ulZkHUPNfxqPfValdltT30Kdi0f
0UNeR21C0Ujxen6JILndca9yji73d+kU/w50BYCioytofb9Bp/GRIKbxfO4YzlZ1
Cq8BIKC/a+4tt/+mS/8RSaAClS0ZKaRiqAZ92VTW/Jv1eUmxC5cgnRRQq+KZpurF
yYohLST9BIkHrpLGGdxnVcfwWnjCFC4K/cTQyQmidZhvFJ1owlfwFAMxFrVRjH3P
iatnGeQB1imFs3oHeWrFML+qqsFAn+QcBJApzFSdOWNnxTXww5EQ4WN2yLR5+Yyk
3NR+lAxvgo1wjSKbVbQ+h5RGq3mGiBKUuexL4hJh2aIRXvm0lF8nMgaF2y+3LcWz
04fOQ1h4C/9x8QmL1a931rmUvNKkCfyvUcVaGwbTv2hnLpGL5n7dHW+oQXGQb3sL
XFhF8qMbK8KEh5V9qJlTgZMqrX6sXW+/MfGZpHIONssOAsz6ZKW1nfhZKNGybvze
K/JBM3FMrhtMejHoex1iCxz6xpF9ErRp5CnExjI0b+NecHK/um0gG2/DTVUBB69B
sX6YzjHdg5aLXIn6jR0gL84HH2lGAjwod043BiZnsEyS+FdkLZtET/Fl3eeObvwf
Aa0r97kC8N5SXVfei54kdjw1LNTkac8Iid0TRNAWxA8qVykT9BTaBXwszXPxsyds
WyZIZ+hEoo3kraU7jGMr/ikSVFwKQmppb5sRZfGtOrwRgjL6ktM7BHVbOXrK1o2a
YhiFY5W+QtFZAHlHsuMiCJXv25GgGjI1x+TAVDsPnhVcnlpAnetw9C7qOG65YNuv
4KQRva0VyERDaXqXzMtU4XNKIfGldFYTD0ommT8ynwh5Jz+hI3+tsE22R/aOlf6V
DurPTON/zZQfav9T+GsnLFTJxphdgQrJUcDDS/4u6Xh4BNd0jWYKxO32zm/2jJpH
3/wNobWFsWW7RkRfzOtW4j+2d8UygKOKqZ7OHdri/RfKMzEsrlPW7MXzRt2QcmIv
oZNETdHMOg+ocpuCzrc17ICac3R8VFaJheb5/LlBj3WPOEnQ139kBnYsgGpohK9H
sxDG/RFqaXxXD97Y+VmU5bfCwWXhAEX4eR89F051SnvzbvWz+svDjk0EowQlNe6C
Qs1VmAUYzMZh5EGAru647g1ospsbyi1gdF8y9VN//q2ABHJLUOt9mtnGd8wPE5uo
yYOIpOD6zd1aG7f8gN2NONjQICWt1DM+PzKHEfjaw+31gvizhSeF93yFVFmrk6yT
QMK97akNnq11097DbM2alURh0LWwKGCLJyWC/ndOIOgDFEfutdplxr7nHpOg86cS
TahL5lalUMLrMleFq6UBJzRLkV6/tv5AmOOlDx65zTBKjTNJ7ypShoV4dhGxyyjw
R8GehQCWvDsUnqppDhfaFM+wpYN2IZDEGuFd0fnE3B9PgD1gjDm+GCXS4rOlb0FC
raewe5tsX3LRHWbWDb2VtHgEOa5NAR2mXfOokn10whyJ81JRqXWe0aEkM443cLhd
A8dC8mfs55NoOD1f1K1fOBKCM47x7bhxm48F2+tl9MOVqVBVXz0AKXU7hK5YbG5L
/2l/RfO2n2G6Mw88NTabUgCWkiTnsheBql9O55ukPkz25vthKyUcy0ZHSYytc/8h
TyGxDXSIe3I8Gbfmgb+e6vS/i3QCPqoNuGmTZ2nsIvKYNWsNXPa74KmZSs7Lrs4O
g/Li7F6YiV05z0olnpeB1XeqhubJw4PrRpgfIbkps9XjMgOKk077xvAfXJSoLGlr
Z2QTqUysHS5GVd4a/okBU+Ppl/pbp9EvRq30W67QduwfPbiF1DeQAItgzL68uqNW
pjdYH0TIJT6MfTsiIP7UPt1nDPcMyWbUhkvra7rWqPtwfE/sk+9rdkJ/USxia2he
TcRlzHeWsbeGIUwRUDJluUqj4lAWE/IW1uF9pUI5DEgXuucJgZt6lkV5NT/Mwkvk
DLoIoEWw0SlI/t9hsL2EWvyWHi8PwluJ5IWZ+A1RCHnbmsLqkv2Bir8A11qlAefC
98/ONEmtPz9BjDLjqHYwn6PIGaEQUJ6NzLxB54Qwan0KJunWtMLl+um1U7CWmsws
CFPQE6gNqtsFcTx6/tY/tbqDCKwq6c+PPSIHu8klUOJgpKdf7wHfH+mGtnm75h0M
L0DNE7Oh9D9M9mE06lcKo4OFiqEhHI+nmYI/i+7Iv8ERc6Fb0WlLrlM9mosa8fyy
1o0I4+HPDFACaqdqygqiALm7KDvwA3Qr5MxRFpKqRPqLg/e66JLbUJ59rd0shUVC
Lb2aGaT0PukyHXyhwYQOxQBOaI75dfmsxJupJM+4Eu35pc5Egb4/7QbTU2sLrG6i
zKjfO3t2stLKdEf8Ll5GnA3ggxAXTeBidW2tYmvpJBdri1g1FaNMx45HU1I0CVv4
KVCTXB8KZu18CCX675KW8qNRZA5zBgBGlIDVcuqkI4mRV8i1hmQL4Q2rjkjErXD+
Xu+ARdcvwof/McwWvXSqpF5WPmD8kh5sdJphLNzS6oKn7zi6iZh454aRkh87UYwe
3tJRTi3sjVGWNJJXnNP9y1OKCxb796hgiOym2s8jxmBQlggwkgzv/+pigPNAGW0u
uFJraKSBV2BCO5RqsIYuFsVR3y8YKTlQk9fcQmGpvPPnllCEMO6B7UYd/MWfWbcL
HY0jj321ooCb4j0Lg+02dTiD4YrzBweEEQL3TQraOSLXuawH9jy321LWxqWMc2H5
dPZKe6uLU7HFk4Ua5f+byKHAMpz6fqHhstarFSmyuJjHYyi/EQzCT4VnjVvHSVKJ
3Q5qC0jbFdqX/pp6zrrbT9wW9hVkJMVckkrdkp9lsozr5WrBvarqDVuXbck/2dL1
phbH45RZlFNnJUNIUaqn0AkdWCcYwvElDaU1wTRRxD5LHfSSFgjDfbZ8VhynST7R
NoWT0o4KXCuQyI7wVI4fOAHepgz4mUZmsJC72dj5px2ew1TSTOsL3MkMpWKqzOfL
Sf6jqiG6qLGgR8QeY9LDmGoYOmZh+UZt07oS2UZ4UoZ/l8Hys9UIFs4SrxHwgrlJ
cwu0Y67K4XpZUzj/BkeuhYXG3OlZmGDN+kDfMNz5TmAO71Uc93oZx8ONEhZaPF+R
IFqudpFjBsenFPdJsNNgmCRvrijnqVrTNP/WamInwwD1/iNiqAD0kCf8RGhkcDJg
T4aICq5bmr10roWQPklxcYeD+07bJfl+zVX3F9Ifu3skJKCbkdr1CBM1bpCqzyJa
yUE96dEw+PcDNx7JeNSSOtMFFEuBhyT/85MMfsFQiapxwx0c/nhSOhceM0Id0F9c
+asidBVdMLCJ4zUX+OxHSqhQLd/cX3GIy+JYj3rKREBJzg1WUueSy+kDK82fxCpO
umFD1jP31wQ477V+6M0IxlJE39od2TpNrVRinbY0BRBq9N4udqMe7eDmDga2w+nJ
GPQa7n8pUJUx1S8OMX+gPLp7QnMHmhGiWqCq4fvD5L0kMZSUs8DMG95JW+xapFuT
2MbAfBgnEEXY4O3P/ryYs+xmEIIS41yBKKLrje9825IB0oD6hXbxUSk75KKrOpH3
P4ciuSPsLoIUgDelLMagF6wmDogLZLjZs4gMU6WbiWllglLg6UeMhCp0ZugeHDUb
Ow9BEbXI53yueZ7MN/aM/qAnXlxKUon+kmjABPBpI1q9AjzEhAkvQRW+Fj8xoPZv
zPwV/UjaLkB4CE5ASmJOJ8HNR/jdTBebepf2083yCUjV6w07fQaQagz9F7eSUL3f
b/NxmZ8/DoJ7GJBheDsDfQmhQS6exrnI/JwYjyvkszp911sGGWL0Ysy33Ae/fSCe
TREOYQxk08X//id3OvhI40xupGuk4zaIZ6Vf9yke91R54gAy6hMRbrqlv1zqnqOb
9p43g0Dd3/mG8xR6Sj+7EAth7pz87nv4Xx1PDlX/F6ui4mONh+RPvVvpMHr+/lUJ
Pq9Vnev9u2VsjQ5apI5PRnMwoD5Yzmel/eyUMRr/P/+mQJ3DhxyBP7TqQEv4aZ8t
pfR7ch662zHPk7z+noz9cV7pXO8M+WE5zHzvDUVAjEc1/JotuD1Dd8/pu96xSr5+
uJwBfLj9e8Tgczvu3V48hqGYcfT+9l/ueROeLQPJejj+gVL8LVjU7GXkboJzh0MH
NuZhbU3iCpv01xEM7rXL0dMYWrb8YowABWLhRzOyWrZqIG+vIDHzCXJ76Z+53FUU
8HC4se58tWrikz8MV/LTEKzGNe03xfSu3Rv+dcq/OuopRVieFQ1cRWCD3RRYHK5c
ATrBNj3k10P9puJAedQD9dC4zE4QS3cCGTJyCyLez01oMJ46Q0cU/2EgWvGnlyCx
bJkUZ0ZE6HNLSoE6jg28z8iooEdkjmNgGnNXSl/6INuy2mLVx5YIjQaKYgtV8DMt
RQlhxAxjUSBECQMgjCjEsCcKibHyAVBUlKCFBF13X2YwKbFYZeaLqclbEICZ0pzx
FdjYlF0HMm5Korn2KIXWsIt6U02orqUSf9Yy5sD4DzytPY/CzvWSmXr03iRIVt2c
SEAiuSDySqlCvsVgqS6+JypYarlNAOLbi30o7NlXuou6Vlvx2hwYN7paHilDEFZQ
Y54fEtQkaupSAp8bPkmoz7tHvWrfIaMCDMnps0+OZ8AT6Oc8eyGp3Ar2gAjIqSpn
ZvfaAb98UlUXXDrn1FxAgTfMGJRscy8CJibUocex5TuiDr4bRgVIWioPq8iZzEUm
AUFxgmg9p6yVN2Y7o/alLv4WHrT6b1HJvTRfcLmGPIgLzq9SyNyd4Zb8jgz4pH1B
eUzWkV2dYgXdxTyN8iStIPhhYZwnqUgmjbtRVZLt8dVpRRQ7bXbDAqqsQ6r0bdkX
cQsK8cnw0mPry0mHN9ezGOxBXcWNy7N+N3YyFaZJ/5TMx58o9GmsxshdlzfJGPRZ
SL3PwaxOZCjdeMpM6hzP215U2Jo6UnQ68DtQsnPX/TuEAGdfLH6DsLH/PFWw9Jho
8gKUncJPX/u5mDaEpehj3KW5i9nOI7NABFPlu8v9/sgJOyqkpGTSuYfqslvwE8VJ
HtP1g58vnMXDNFWvLgMODG7l8crA3bb6DJTnYYBc0c0r7w/2xcauB0l3hd8ZZGaZ
u5M9nUNqafGKSJMA7zox8OxseaT8tlDrRJHSKrhch2OXHNP1Fy65Cw+Pzsdhm/Fp
wKNyttIdWXVvMQh/cq33+befpZtab6eDUHIEynSIdedfLG08GvHrTMCBDG3R61M9
YQpP3nnZ/E/zqF973FJpw38k+3qD/mEmkmPqWyAfeaHN+mKcximx/dlhNVoqaRmi
tDdLCzt7X0Gfy1UEFHCKOk0XmpHKPHa5NGmi/Or8wY221YxOwyIFB4R/lV16eM+u
0qZuLwHuiFSuhbUQL5XyBxjiaZjs2UAbY6MvDi3VsrYnIf6gYlCgMBMiAjVJwxz9
K5DRRqD1i0NWJI7+LRAKRBdmvPC0tBr5AA2lo9MyOMzL/aDICI438/fsmetCslvF
uTsVKODLGrxvaOH3d+BTuTr496udZ8pVBdqkR2hjYUqF8gY1zMKUXMH+uvekYrc7
QzjYbjMX9ViRT+VYqdUnhVrLfdtu4AoxoJf3jLgRYX3y0OsCVXfSBj2M9hxSRquU
u9IhwDtxLlmvt35R9IFYtSV7ElK8+mHtzo4tSgxpXcrS6DcyfAcdkZ3UNeJxXlYv
xM6Hw8x0Gx/wrcj7TOOkxn7pEAtUnUxIW3kcTy/3Shj/Z/VoonJeRBZujsKLWNqX
WdLrsr8HpLk5mJO3a/bgq9lRrMuItHO3yw0LQjUETStr8BTz3skJ3sNeW1Ju4U6c
dcsQntraJOe6qNdM+XAmJPkmLph2/LICvcO+2mpXpQU48rZsQN15fnds5UFAwXVB
Key3ndLX0EHMSQiqTx8///3EKepYG/wTq04XaIYo8QTtilW3yHQhdpdTS/9+EwB0
1bXrh+hX42VQaab7qT6cwuyYP3s2lcSXhn4Rvak9Kw0g3y7Uz1UDukm9UVHtpYc9
8pDZL6/fMRTjJwEiruvbNNYCgs6tp1NG+JiB6jz725fsaP/gFzNQn9lkysWzl1iO
XBNTDTaT/KrJsNzstVNYYtwcWI30hhfgW0jYJ7tKmPcWz43yRPRDa0UV/zSyUF6T
uN4FMqlaaFX/x7TcAVr6+etw+n//9iz8T+Ri38Hi1c9eAEoP6Ag+8BOFCMX9/EUt
oC2DDDOHedfP1sAJAJ94hj1lUrgGbqVqZYduHrgxhKDgBwev9m+RgX5T2BB9KsI/
98NFMO7KvgQuyt6rcdSRrus5//wiBMS8U5b+ZHh1HEDbdj1TZ38crtH/fSDd07y5
10xWjsiSh0+JNiIZl3IJdEpl2H6YyrBVMftCF30xUzkFrVEuMYP+RdeWMX3Xx3I1
WTic8ToV6mTOqTdT052VqbvgYwziH5LWa62XN5OdFpY69RAcz+4GRGYy9nxCoCTF
reMh8/EuRmyvkND9aumZoVJBVwx2nDDoHVMRiRktsMkllI2sn+EDOZsLaV6K2AE0
4P6idEhZRtqOvZQyrqpa7wQUBhOPvWKrvVbpKp0Z/XMOaXxwVGt2wijOpxE8E40g
XdEzU6Dd9y6ShRSuO8ELDZxwOLk1yvt3OTK0vL8jDAbqiaenbpvpN0UQTO/AEtD9
iNtk+CZKjOYDpje92YVBhlWF8NiS8O9s7aWL0SVjFYdRVxdt+Ccn9eG9iFaS07iE
rWSPh7HEqF3sJalz3zLjtN9iiarpqgj7pC2G7TqNYQzwTYOR3f5XlbywVTxyMCtA
HhFtFICTfPLKYHlkaMW+2zN4Ngb5idOScO2zr7VXyIBxt1hErI8ghVA1pLdId3vT
inJhFOVKZHFnNVOmX39EtKfLyAVkJ/eqrkRb8CmJdNzWfulaTJRkBOpv77zAwSVl
vvFcFaZWrsjSUu75Msud2UMya246nfgibPhpme7xuydODX6e6PNpFWkdS4Pa3u0u
sxS0/omYOkD5KlNQeZpOu+6X1E98UGC4Ik6ivsp28Ul0RbPRx+IS8GsNod8LjjfI
QwQ225u+lzZt2st+hhRtAExOVdaiui5zmtXWHhKzOBiDa8N+kfBZcwbW1Suez8EF
BnGwV/VxNZ4I+EUY+H3tkxnj0TJ0zfd4rGoK6FQVJ98cKBroxgppVG9QTXgQI/fZ
o1vhXZKFQeKRK5xn+XrlfHQ+fEehO08UvPRVW5okiJTSw4Qj8AaXbod7Phxn9/1G
RvzrzC6jlvk4TGHFLt9yADBwqYYJ76g74W1SRScyM6h7esALLTGg++0wz6EsjlKo
Lzt+zfR91lj05w9KXkDkknRTRt9K9mzZiHRaFkLvD00Z3VRVE0C6Acb1gf3En5nM
/tPASwzVrqSRo44oqPu1E9GFhnHJQ2bOVBOagxmi/0w2g+K77iKjKkgphOdn0+4X
tT7MYWktMG0dMHJNVqk9y4uaqotPaWA50tzNwKXNLb1ZoqlL3jIBnymDF8ijdPDM
bMSK107eXXX6OWWXa38nGDtkmOer8DXyU2vUhjtC6OVX5CZPNPvEUPoBxYvkFkqS
WkhV/OzmK359R4g2amT0pDfe/i6XrMy1iyBClfy34xzdF10NsXExj1FlqKfnY/39
5Oekojh+V/pLiAZOQKgrtYdjf4ADFdwfGhnkwhPj+vE6PD3Dof3gcOw06DBOWdQG
1/VGqyMJ+wTngcJaiq5hdsF8P8YU0p1kzNfa0RQYiGH6B6ziJB/bLshz95qytkax
zm9bb3UDumkb3p5Vu/MXH8JOuuMNZSNgwaa6OaUVtQ9PLNaPXoQ6tyasvIgWXLcj
/4GRw+Qc8WWEg7wD9WsBazu86X1Ov0bnBjIirmVKa3QJjuP/PSAqHMqpZmcl5CO3
9ofsbJpqEsonbnEi4vrhnmZQlTicgfsE97l6oumT4GxUMd8yGZAe7LIp+5dRm6Om
QIAtK0QRnmVOaS5G5DKORI/mejHIBfYCLBFxSc+2zck2XJjWz3MyCTZBh19Td6lj
bb1FEh633uJBXKnIJAtubihpkIt8YS6gTn3cJT+4EKZs1rk/nn01i1vOVjR2uwCu
WCGQFkfLIyZFwkHI67IYYAlYKFehauaRTTu+XwXdnw8WRr4x3o1hfNj0J9FzjdIH
8qAJgCJCfvjMZm7720nV432ERBlbJ4NmmlXKpClHzCtWKHdPzObyNsmI1Jy0mZDl
MJSzQ9FR3VL0ZN4gq/D45Ys6/TMJD7ZVHUTDLUXkWEX+Y9DFYxWkZu7pX2gQwIVz
uEx/QR4wTHxljjLrM4ndumF2DBvJt3QJsnx/5fIdDotCE2QOVPhAwmpohcvkcrzy
imvgYXA1YXVPtbMX+Bh3ShF8kWYOZHEs+yioaatlvOTCx1xo2lIDHCXhi57BYRXG
xjE2NqeyY477LLgqYGUDbLtjR7SbjfWCZxxeRKwMyBhR5WcImrohAoyqFPQCWgZo
qOlvZoVUuggYfxoA9BFgo9qEOv7G5Cy7Op2IDBWRVf0r2dD57dT0AztwO//roi7l
+5XsTxd+AKJt5V62AXM36XuX4XJZcezBAAK2M5EyUxmVi+SN7W6z3RYYaaM73wQd
4nLbcbxJcuWMJjD6IxC9T9zrHppbXRqmtv6arXNcSfsf2uUZ9kApAWFg4QFXNZU7
su1jHXMlWEbZkpR6EbJXjrl89KKQS4Fvc9mmWFzgThWJSM/yKI90L+ND0Hc4nk7R
L2WTboFQz2Jp//4tb6fSOE2WIB0yI36WCcz8NyK7gveawK6jDKvLQ3N2uRrFh3XX
ea7ppKxojQps3nzqY+h3e1Ho0I4vJ4dUuA5Z6La2b3VbwvWBcTTUPS6AY4Z2tbp4
vQp840HxxovN3QzKAtvZOxoTBcmoo8Ki51+sycQNNHrbNxugVtR1YGK3GEu2Ljjx
z+U6BocEGo8iuhXfLo8MLTAraaO+5v99FRbq2uvownTV0kpkIRKbn8EixGSd7iIB
LN+mYv80J75kS9PBa6ZIURC4hMaLL5mHcBSrNtwL33g04fh2VfGpEth8qEEE4v6H
KBCv6OQ5W5YBYEFaATs3q+8drS7dV0ljfBq/GWozWV0p29uUZAkQW2USsRVIhmbx
UCoDZr/Ax8CheLNEXoup+jKBfIaTyWWFpeclN6kj/nvDElUWxFoo1W2tSGHj28tb
8dBuDRaWLx/SQOuySWPqZDi+xaWsmyOlvaZYPtDLj/KF2oX9Vxatohv7qklPUsnP
9fDTwEPqKUmoQZolJR57S9nwpaTUA1Jpn9aBgd6+2qNtrHh87KoFGYoO5BRExaV9
XsHlbTaW+orHnH+fq2IuQLAg5SRS5ju6gZgsMQlrH1cFCD0OT9W+YodygGy3u8ew
VW+57PS+Of13JD57qkTLiB+EE/fNaDqQ2O/0/CFKELQVte0bFFdlxHPkOR31hsiX
R5gxq8hVzq+8/x0YFqQ/b1+9vgV56RfTGwPrOsQUOYCIDO81t7Ca4nfvdSBi4nAY
pqUbs1Uu/Y/xHbCQOP3FIq82zPN+Mfn3uwh5s6fgsHHXAF+uhGMb0muepVuLPAJG
0uusGP5sER0iF6sI/UGdHBdhKBVOod4twAIEn37eVZ4sIFL+GbcJjGjO5ebIldgE
6NGEGFIcP0mOHSnA50XPt3EiRYXVKn4+pWsvDY+Mku+uBvQY7PFJGa3i6dk64o0f
pzf/HEWshLvGi1mAcPqDr0cmogy3jn0XYJfSa+rUa0MeG/yaTjmw+2Dp1rksUUbd
nhaSnMYMyfBCXaMgTIk5wqXVxxZSvPkG6ZrzwaNqnrdL3UOPB31JY9oGS32u5gNe
1DW4KH/QfY/3FhPhpV/5pAuoWywbtPei6AwqLLKXgvHgKCm6fplo5R+Nb/c2AAL2
/uhkcUQ9k13wlfjoE8tkd/n0IF9DnSlT0WY/Cu7almRt7jWVHKGiNkECY5KXrXPU
ht4m0No2NVmiCtiLvBm/2phwYcPRVxsXH8Pr5QwGqMCJ9HSo2uM3fEBHwaX3JKGR
E9jaHkzXbxqfRwXKsaZOZgkMCzGee4cYP06CC0lipk1U+l5eh2L3SYF7PPgc7Dlx
rmNS3Oj6Cj4XAqjbMTbFGrt3ZJb79QS1LqC4OBCT13ijYkmyBmt+Vo7clh1nZaQE
vITpFnECMsg6gviyXlR3b57Ag50na7Cai09HaWYldeuUF7sDi/73GCG+8HjeSLBM
pblXDlXAA8+UtSC93RSGo58+GOwTOOt1Lc3gEx0MjR38gWcLdlxyH66+3CT93WsL
nSBmgUN1jxPTN6kAFGsYWiqpvn393PJYVLttHPQukp9SSPSt06pdN/BSZT189vp8
J3zbhb2Vzy1/wN9EDJMR1/Hpe+TS0C7rYYoZWxIRvGvgedInUKMbZCdm8TTX2ZN0
EeCr6NaPCOSnVb/X5GlwFUVqK/wqrRpiHWMD1l5tSy9ysYpwGZlv8h+onB0fYHnQ
ywkxCsHr6TIhP2mY9r1Mc/5vrqsNy8s7EDyQCmwqgcuwoLdCAFvgZ6jKHVUhBRwo
gS4DjNP0Y+wAaRWPmA9FTkalf7G8926ez6brsyMDlYFGnFuotDzUSbxlXvXRmDJu
qPIoWg3Y3K/za1Vkkdb20eNsD4/wGWrc0ap4zX6U1kZ6mqiBb8NqQ7rdtvo7NY5k
spCMXoLaPvS676DngC81dwvFe1FNqhvi1Cqlmu/ZePx12P6CZrbTcs3zPOuAtrtH
2/P96Gt0nlGqxoxpieFKj2svPvP+Rp0g04beuPxhKhdsslQ/EfaHfcJRMwSHeagZ
SsSJgh0XNRzlNukqGvpMqS0qW2Di4lGG6Ske4cY/OIO+3OTKDUW55hwt+BOGYmwZ
vEUX47qLzmxnocpsCbbLNXywcveWVSHyFluSibgCyVnvMU0f4uo0TwoStCGWBa5t
rMk/6vPh07IPFrwTn2Bkh+9Iy9cpFz4ceSWNkAXRIgti+yYrmo9mLOUPTSOOgxDJ
JqqxPIpoeXs2oPGF5pPBQxKSBBIDjQwLqtzMWm8CXKUZOPWMLSVkI86zPRpj6Q1J
dqJiCjKbEqXGjXM5CoK7boyIJgwja3QcLFzsKtKnRAxTtyjJ2x1YzqhR8F6obtf1
tJ/jhwl9CNuJVbh1VCFFH0P5AQ7xn29L/lve/V2BLCgsCvol9k3Z/t7erNClvLRu
5E+jy0dx1ZxHTqnsk8TllaJVwDZTNZKv3+4OHQwgjWMOGXRMfzqoB9ODJgAaeOWp
b8c+P3odXl8XibJkJeCeupumHejL2jRtAoAUsUvcQKVnEi/J3Zer/AootmSJeA+9
HLtHzZq5MfKCBiJHYPtpzO2K0aMAO2SZVR9rjWJ5q//GV8cszrzO6i5w3R37vLrS
P7hFwKvVk8TiOXNMsNm5/pplA9HMso0AaaUu8Ar914pZBDZb6ac7TPxl0fWRaPOK
uiH01xdUYpJNWToY1eFqhm7uZQeDkY94FgVdSo8BwVkeSU9rKyQsujWMFFYDaxtH
8V2MuXz7BncdAJeg4Oth7BiiahMAeEF/b3/V4SkQ8CXLaw/iZz1YRPlxh29IzHvp
nI+wh3aHZ7+R+dWafL+XiZ1JMQQaJdADgV7VENDcfRX2w1TwLEVe4O+H2ghPooWA
X17YfaJvIZWsQrmX4ze9qoGesj8gzuCNQdt521PmpIHVnIVqS6EUrOUrkSHAxHYm
goEEfQkY5FCjBRmMGKD/q6eebqn6d/C3v56Jp2BIIShi8DOa9Jfpf27CuXv2ESjF
lQqh3XaS61JujIMe4PONQNoq0giK13QuvcGRyA8sFQ7csevqY8z7lHu+n7roc/kH
GzmZNHC/kQg2D6nprzHs3NaXnGVMHGIySk79GH0THDPWw2E2pnpb6Sx3UVMa2miv
GRIEmdAhU6rOU0FkOKxX7qHIkEkTiT3oA0OfuNSooi0IIdsMZEt+Yh36LW27nL4k
9EkOXFQ+ZIKwBSitEgfutpy+6p4zxzS215BZevAh24oI2+hCdnGxRWYuL91S8F+j
KshWOqfwdLuKrKarpi/kWnn18JP3PzLnJ7Ada1pyZNL7uq5onjtzFcnnIoNucBaH
zgJKPVXbdSx+mqKAMJ1Seq/mmXti2oSzlssxMQztjNfbjpfqj83mSxb7Vz6ESYYk
wzf/tITxcjK4Hngi0Qo4rIGCfGqDxY0vOOrLHAMtATgBBK6FPickDCJ0JHW0gSMu
dc7cypqkpeU26CIAH0jiLxrrNB5ZVOdbAZom2Sne4T+Je/X5KePkAC3s2sHueuVJ
jYSxEnj2bViD7wo4C+6dRpkCMKzWe4dqqWz/F4CudaM0+xJjrzgxxGw0Egb5+9OJ
yfAgiDAYABSvJW6lJrCbDJi28mfBnJIjtwzo9VfFdlOuX2oX1nGPhOh7eiy37CaR
T5gRunZqwTqajoll17vYdpz15vrWJHIy2a5sMgdRZPSfV2EoIMDtikXoF0rwHcH5
o3Gf/hjlUdxjNMQp3oIgGIsOhgm9+ghPFihY5sf1Esr6J5255kgXV/nDgSlEz4O5
Bjms+5VLpDqv2hG9pLM0jwE2TMajfQIsGhF3QBrlAkiMblCXL8iKIi5M3Zf8qoFH
Nd0GyQofJZSFvUjpD0gn/8QL8yXLH2KpIv6tyIsObrIqq9esUD1Mbtg6ve6UU5Xb
i4VNu8ArQcqkiH4OBXG9Fa35JCZCRDBBO+qVTrmu0vbY1wDj1CxI7RoJC+CRPsmD
LP7NIYSPICm43iIhOBT667FxsBQVtlcULoEhVLtc6nQ33vnMdHR7d0ie8HnBobuY
6z+lwzZOoD8hCL13en1NvehVHLmyFrXVggIlASt3LrCfQ+s7aBxmJ6GGU0Ay3TSm
em8W9JyLuBHqEIeu2qUJY99TsfJzD+ld2OqIuvh2lh/WsFqeL2rVqTNA03p9kwaX
G/xzF7Vzr+LIhP4QbnpvRYLwyFYEFOS5lfskZTDYPt7I5eTaxGtPPTm89/3sBKyc
SR77cssEMp4cx4NRM1QMKNz73BJaR0XKFyD7b++zB+6FqsUhdBrvZLC3iiY3qKmi
7l+xpGp0VjgOHq1RoAe/4LwXe+CMe219GsVkhwznuz1Dq8e13Gw1uHMl9TqOhrsl
463P+UQWRUo6vSCx8FduQO+ZBZNreplYSbgRwAmRTGsraumeOH+94ViP9/tmEay+
C26bVfktfkvz8JHIV4SKUeaBnFxryM5X3/kuhGJq9ZN78feyZWO1K+3gu5FCj7w+
0Tqv5n8ln08ZCFeAB0Txl2KuLldCM+PKBACJWohxBeslq4A0LalliQncSGOk1sEx
G6ojSWhEI1ubcfjRqj/i8Fbs7fmPQD+IFJd7eSznPRNMvnS8i46TBwLVK4N1rW2R
FDJlzmH9qQOPxm/tJtGkASl/FteuzzY6NzT3gLYBKRqFuNMF03EKpX0oX5g8AhlQ
oaCikfMytK2qvtFTjNgKuTvkm53/SRwOc7CpbdBCsu3wk2cqBhP9b5d1xeYEP5qX
DGikA+IEfKk38j7RfNlF8h8g81zyuetJmeJpFJZ92hkd7GuzuGHBpBElz6Wa8Ow9
+IDbFB7YgFm/g5ic8/Xs0/alVKkC7N2i6XDhMzHJIipKibD/0bJWg+CtN9t6nDMW
vUQAM6j8w6zV64mYFmrFGDFRXaW7lSDSQlWii7po24A4jKWpcXwv+oVm8d2K9Z+M
U3oguHbXVUUgA5noEm3USk1P6y/k7zpr/NIpzCrVvPpIHGZ11oo1zz0PKwrMVjaM
1IPbXB6HpNj0k1BVL8ZzQyLYNpugDBHkMG72O3dR54NqpTHjvC+wt8Rln7PNgzyO
wX5tQiP2Rv9hH7K/g+j7pwC+ucOUhAsJdhmdwsWdlYBgm9GVM/yRMgFzOz7MQokh
FJoGHSNiuJ37c2rsrru6luz3RSzK2WE0j9lgpSazCkOK5K880gfKvjOvFW3PTTvx
cHf/OTO5Gb36zTDGMxKtDXY/l83jK+opn6b4j0txTUkzQkBmls8nb3G3Idd/dXqJ
FyBBYk2JuX7Xas5w9i9ivw44p6049/AceUdFexyeEFQ7YxgOupdHTcTxYm8ybeDW
D5Jyu1VMsc3LTOJ5PbJ4fbOlUuWc+dVv/VyLQpnG92ND9mwVB4w9FD5QDb6XkVbK
ATlGgozP4pWwpe+3ixwL0VBSG+EWxre/HLf84DwIV5c21FtPvq6hXa+YIY9MhKdr
YZmiHgZRS/V4AXt6dpAZ6iHyZHBuB/elf3H4ezLMIwa0HhrhGMx2DDmcnOMbyXfO
oUk5amveEC/hLB36yoD+ZL2vZTZ9fNkT2789/Oe/uOXyJco6rR9z2Xxlt9vb8dDQ
r0HUjitezL1KI4PeTk98oUTFk//u355QUDXPfRYMZ02Y6ldocmig98dicyQmGumK
mZgvmYNYxJX7Ncu0UVqEIZp645zlMzmCTDdkz4k3A8EoG/m8DmgIBe6yfFYoYvOt
50dabcG8JlQma7gdSlDT1Id2QvvNfcgky7ExHmEYoehujRa6M0VkGVTLxNSj0N18
vezsXbdZEITsiTts6HH3TauaijwIyKvPAAmc0EnyP87YiabLejiizGsXcEvb10Vg
4eZiQowZC2WZpYZd/nFoSO+5KTsSs6TYmO7KIYaZzBaZMZzsRXN4J3npBO2D5rVB
NE5i/a9VqjmQzPOBplDkZTieNikNaPxuxzXZDQYqyXCqcKZaYBHt+CCDOxjAMi3o
R2XKAJxMmaLJv91BCLk20vQQXj7QmDXgChQwv8vjSosuXxr+iZnFCv3dshmMR1L6
DaqAgnTXqxrlrxmND0Qaz/dip86uaBngIXk2G3GCYknQSrmoJNgYhbUgzXQ0CUBz
PHxXbq7ENregyftVxwkWdkyUA7Md0BYp5CS4ELgooW4Dp0oC7Ay5uqeAYOxremur
ZgtkFzjPBPfGz9Diqt+WBKAeL2k2LamJnFRE3K2h1QGmvnMLuw1m+TgU1xVRudW6
Wdk1COlo8UDToAPxAnvlXmmRvSotk0fvRgM8Dwgt2IjTdCIoYc03noRzs1k8+bfi
W/b5s63vDlnXupsxxnpmVUjvcYcUc4lK79H0cNPQUd/WeqkpOpGRk0lLtCDBCwOc
DpqGOkMGsp3UOfVRq9/OGMpJPL8nnXWI6eO7/aeqUl05lhbqPWLpJ4+ayRqSnXyk
M6kRft43btoUHYvBy5fN8I9XEa3suNiSRwzFl2oEhDttLEgMk1xJpHEl+aQ+UMg1
6XlOHowbRDr6XPA2OfUs2c31Br4uwD9OjTp72T6IAN2b5H8ulq7PBU+vS2ntO1KA
CSu5+IcLKszP5RQ0zbMTOZiORLW1IKwFK24pCJqh073g0NEJ6cRgBMUgi12s+oci
XIGMu8fjjhpvU+G18nC4GfRaXO0rZbdgWOijKQSIzonr5pEvzetSsq+7vuorUyDC
0ebRrjcxk+QvjMs0tEsJvkE4OB6fm1V0UUVGhym3ZMybOaE/SufR9MshjOMYzNRf
zXTjesHdSFjtHsfsI0hM+M9yaJRPI8fCwzl+8EhvgXtu09YUGEoiMnQy8ZYqxrgZ
aTrQEJUlEN4haiF43Vj5CdV9oV+vvq+AArgp5USc7UgqG9sLQ7VK9acEpZOwW5eA
ZfRtbNhBDO/3ROwhasToVSzwHU9WC1zqR6s2kC/iAE+nN4ZyR9T5X+gi1nLBxEqE
952uVVEKAInpcrQ872JoSELeL5ZvMu1bjH07Jv+i15pahtWPCX/JkkQ0OGS0rqCj
Ydsqdpp4ifP5L0mn5hcguF9//Gl4OVLOCHA8rKqCufH0lxINZNb9eXRSbWxnf18d
fQQxH7qdG0q9Nq0ykjp2ugnjWIO3R/NAKlqh+VUTNGUMoxcQ8FShNGfDDn2n+75l
JFsuVg2g98s/kI20migv+uyd/Mv8157f4D+HkKKMpeCYNffewanuP6B9fOBVuG2v
cmWQ6vbzRZq7i/YyjN2PeZkJtG334LDCS2u3Mffzh5opEdJTGaQlFStnGIBl6GDX
1FlxYQnhyY7oU7gilJk84cE4iUTvc+pZO9rk1/Xp6UCwaznaFu78PhLYX/c9rnNX
n8b+JhEdDESkseKQM44ixodnO9oJvL6aPDw7fsYyjPw2tICLXo7O0cRbxCmeDz49
J5jG5LVtKMzBhoJxQoZsEMQMKt6G9nZ39TxR1E4Yftkxa3ojUYjWRHAnBgYip4mS
Ke8P4ZT71nmUOIg8jdvHP+d0AYqwX5YucwQNksD4LhINoePHv9eD0UTBXqpbNRtm
CkcwwHQ8YRr96KJl5F/4tpAEYidhmNGHDbvNKZrZoufZHv3K5/Fqn4AGld4f/JzK
/k8WV+ZHHqv5c+o0V1POTovPVLxhHvbH+nmpde/cstGAzW+InXpbidGnBZMi4vqu
7Oh9Adi71zXrL7PtTbinpiGOYVBVe3xopQXqFu0quNl/pbllGE2QR/Xm+glOMOSX
Xe1FaGtW7w/vSKVvnf5MRk0SAdv9tZfzS87FPXoXGSauvMTRq5lDHgDnm/AxQmRH
YkHjFxLApV9L49AlO/u4UWrL5L+R2E+aoVjKVwF+B1prnwA9sxw89vwQ+9dTmDTO
dXcS/gT5LlWi7JllsNstD5ntJGDUMHioBgCoAsabtCln5VUGJCZwJYpQRLLqTuzS
PfSbqDTpctprD2lTOk6lKIThWy4rBRMAVVelT/qg3rAQMRqTsZ/R4FP1U+N7aVKW
6SZYkUWTVi+b9eYMbFB3Ur1j/CKPiLLuvv463UcC3x+TZwsG2znlsMHpES4W0N3T
5eFPoNgJsVnwxdgRXR69IdaLSroPUctYQlaRVo7bwDINebB37PJmWy5yoLjNJDWO
WMC3/sfpW+/Qd3g46cq3IpuJJmOpsxREhykw6+CVwittIqFNeTyZi7KFLvJ9Sc8B
XOkF/BORt5mLOlsH8/HJDdPjXrwrV3FKbyefHV+wHXlK4/NKMndaiMuW4esTXMcI
60vTPbDpYd9bGXqNmWOrUj3la6Qilx9GD/8aS4DNTm8hsUdgR43eLAtEfJGwSXtm
sS6MJrY3ULmg06Qte81Z8TGQ5mA6WMyHelAZE2MPzSG4cAPYbI4X12B7w8srKoe4
0lXiN9j+NGB6GngcGz+HGpvxE5rMXk9mGiS0EZutpFNMWu0Q7tPJODSJN+7HxWbO
KuBM+kbyc1GleBp0rFSPOZ3+87Ha3NAv9NHuFrp/wcOOro4Gikv9/DZnYfNdA8Ow
o8cqs8n8i2GnfbGwTi+KWcEhpicbDOY+70I0KAW9FjYKM+NQfzsjG75RZF3FZMBD
Gf1aQgTCG8WdvMdqACSZ59jBAQJM74oRwypXYjjXGHc+s3hdrLDl2MiZidBkcKIc
eivS+d2vDgNaMFfvA28rbmKs0HGTgsQ+snFXFaA7UU40WAIiJkOzB8H3SpGyLkhR
ckuJlG3crn+LZ5D2pvFpZXJIotOwXNMi2UODP9HaTcB9Zj0p52aHe6ByXX68dYzh
HQjekiQduB0uSm10BOv0GJKv03OBupER1JUKRLkaKyksLUE/+G8h5VhOsQn4RPkM
cFgf4D994JsQ/TKLAUvzvECd+fPNPEVNQ9NXZp1QblKRXlIZwM+RUnpFE8hmdgVw
DZY7ZpXpO08Bp806+UH53yFqU2p+XLZmuOkelhg9tzUfIa36vYFUEodT7hf8bnpq
f9GDHrdDnBFxDAkPebcdKYzlGRxPeQg/84p5Bn0CclGiUeE/kkhYi6OwmVnmgnQW
O/vKcyWGm1VN7JDUBQpcrgXs3o64FQkf6AjXg4Fc9a5oes1xfGqZs7xL4WdZFPQb
bTftMy2CRHWFbfLBnEqlNXkH33DB7pw7893ngfm1kV0dsyClbuU72q88GPPFTIc6
ur3wrOWDck8t0F1azf6PAUsvhyHhBIB/uPcMxXwMjRgSl1hIYcsc1+o9nRPfGoil
pVSzfZ1TQRdLZSx5r5HrJ3K/Jb36PmO8SmYcWSThmgoCZ4lswfcDP6Akz3CWZp7C
y0jbAYpvJ0gvApUggNLXWGknEFVKE+NeLdtjQJzAUQ6PeZwtW5kkfj6BUiXTAwbz
XofIAQPyWw2hFT6iHuWdNUCSQRtwc5oGslOGH4ceGaRVjYXOXwgc8CGAGL6uOHQf
cOExfMtv5SDsgFU0lWnbQVACfACHO8HbLds5hanvCmum6chGctJxft+u1lgavASf
e7xagmOOPC/ye7BVgCAvfOIw0YInWvgUjvXtHJljLo7KYamb0PDhxyrxYYb/FGzV
NKlPjmLViHe4xDDKKyklfp9cxm8ELXoYKZkFyNhvLlu49LLh/nCHiLEhOjusk/va
0sG8qXUMa/7VqIeN7EncftGwOIO/VwSf66ZzU9mINYD5k4fno9c3MVlyhSeRmlfg
0Jnno6agxnX1X33vDFVDyNBY9NGk8xDwKGkYEcnlyOBbjDsSTmnDEl6/evJ0h4ux
WMOya4edbRGBzYDMVkkB5gCxbdFWNhS4ZI5Lbtn7vIhDh0MgCK2JjUAa03PdaZxB
DOAzYQlfQSqnm1yfH2bIl6giLg6zgZJcN6/veyX5x/7XBXCqNMo2ccQLv19o7YLS
cQzS+m7SugWc35z7Lc4ST5/4jvuuwHAwXgX9u2XPqwZzzHF587VuyqC8uE3Wa2Tz
EA+ZQJS+Mpp+L11ZYgQx/rsvGbB/WYRUEutmLaCLMWwEUJZp5DCTGQrmcs2KUpUG
853J2nh5WWySijVmqXhNIV6aqyM0S1SG82AtNE+yLwNs9qGCnFfnL9hwaaE7xqqR
PgiZlqThhBfi3Z7ZxlwkbWIgiPt8Xj2sAzn5nM6PQEH//mrT2j0cha2j+CgqVFii
OPbgewGzuQq6h49Pkx0KiRqWnNn5FA2n69pY1hDGRqP93yVigSKS/kKuojL6vRvd
iskuNBelL+mC60VjS6oldvmC3nc5MbCCycMzF/112b0VPoEIg2jvlTf312jwOZ2c
dGcb6/7E0CxQyWxOxSLAnheSFzpeVKux5KteQeM9ghiIMzs1tm3hPYqnUCZbNyR5
8LSWDIKydwl0GOI+RZROM6bHLoF/dVVwVSNdB+laD8AoSKmONCM/uIt23N52W/sl
8jS+Tk7wszl5XOyPIKUJOUcXWPraW0Uorj8jQVt94YsZjYIehiJVljo5OwLzhFA/
b2wiWpEMJxFMJQbj+9Iy7CRKQO+WaCdym9XkoPkusIGlG1hRMyVm1uDDDbo/K34j
vsonx2S1Hk+XC7kvA3WgL8Zx80Fl/ETJXME9SMNr19GcCg57eb11P4O/dTOZCYLq
N/zpaUWNWvmRV51FAnBvp1G4hqBUbFaKjcOtUn6KvJt2fEPkqM+P5fIQli3o5PlM
8G1SmCM3ZCD7ByEpBX4OrFohgt7bf+KOapmR1zTjaFOo/rj5yJ+3xChN890i648a
ZqNCcIwuY26C+3eqIjSGg/oiAXiDX/MWP/+UAn3Fg9FIj+qAU16MgRO8ddt1bbcd
wQJtzrpatgMX7ByxtbKJoVWbmlYsInTiQCV5E3zS8ReuFDRwvtD8xfvvzJr44CsM
mJDJXVLHB+k/e8BH2561AfM4hUOVmOIdw8YQP8IFO3XwIq7NgNybIphOwo6tDyb9
KRQN/KA2p08NV8PsMTbEP81E/1ZejJLwDnjIdsHi5FlOP5CkzE5VRkHswLhjWMS9
oRzlVVo1LQgVdl9TksUmqUznpYuVouJJ3pWQUKLZB23xv8yW1McyU0mdc7JfwHLR
+neaqJnV2CF32H/ZoA9+Bsq+/XiTxgGq6Pw8WEgckAFs0Upq70GK8bylFIJYLShO
KIU01Rys0u+lvDZujLUIuV6bdUncGFE2qWdizEaXZep+BZ9Xx72D1KeTwT5DYANB
yfPX7npvngsoOWhEcukaNtGMn8kKgCXxSi/EDwe2QoEpKaOP75hfGKgDWMz0ZDtR
4fr72vNz5ktuMnk8RrtKtJY+jWHxcbrlN45X/cSPk39yWVMiGP35hOP2DlxWEZYn
KsGJmmwtDm3FvYNK1S2Y0v18X+Ucpfep+eFEJL8a+yuhN+jlvCFWbG8ejsvB/fOF
r20b+sG4lVTfZBJrf4AYkYGwNzNVaZjDnEQB4Odgi4u8e8hhWzB/dPRoSERvF00W
HdUir6Xq6KvBf5shKvwTfnMIeMEFm+9Dh1bPQ1mHG81TSxl7Zm0wykWwEDy9EqYJ
Sce4hbiiou7JUTXr2FUN2CvB1JmKZIqlaK+LLlmLgXvc7y2cn1fYzwkm3Vm2YkFK
1CVRXSyr2kI29rKFIpKj7/RqiNl+pBP4VSwPqfIMUrxywcr92JQWSdkAsXe6DhqC
0wFU5pE0509g4hyA+6HnRmPrWw/8NmogpHfuf+jmfLD6ZpGEGb52NMBpW47172N/
6K2Kl3/XkrWeW1k+pHQf55ZeSE6yRlC8IGDazbGyX4jJkRKegoNYGvWCPLsB8mOX
LuWt1vkD6P2VeRt/OrhQqjz48xRiaRsaQ7jMKUlSAUAPNx0uBu5mkMU+MDNRFq6H
8n/nzaPeQe1XdWnbdem7rge/03zImqzlUN/i/fv/e3DLK2PxHMoX6VJoQQwdaQlM
o5p3s0F5BtuSCmbj8WtzooWzRRpnA6unprdryrH1u9GZPRtiZMZVYt9JkXiiEp2s
ClcmetyXAncZCx0YXjumOiuYAZivdc204oR0io84tj1V20f6G2tVMW9bGr5xxpBX
boNxpFjAN24QRPZRSba7gzpPUcVvJUvsv1SkoSzDsKoR8bQnylJMshHveAHRP10I
nLKjPyp6Fi4+LxDL/p/CPO5OoUNyhjDBcxiyRg7PIP52kE/k2BFhOR408Kb3MCbi
E88BwwFji0n2p8VajeQEiWQByeEijy8fhCTSZgFGRTsYaC+1JhJG15BIGz3Y1e2Z
/oD5iJ8s7SIKY7mItSkAv5vxwJjzTfmkFpNSIWCLHXNwLK3xVrZQzMXSPanRkzsZ
Gi9hYtfGTpEa1aBAISvHWId0pH+s2/KWFIp9Jvd7Wn3AX+tzRTOgPx6xdwIYv/6r
VGdSpKxdTf6f5BbB2YSMdpAUTPCM5nuPjYSgw5S+X4VHjj1nR2+mx8b/J9xks5po
w+RadN7dc9VlUCBuk5NM4dkJeuvokoeEyL9fOa//of/Nj5wqnbT/FyVEHkZenEvF
xJaaGrowxkmGOWDIYKcnXEZ3CQ+NVyxFtGK1XytISN4DmX3Xpnp9J+ueAw+Mu0JZ
c/avascVN8zLxQMlqQXE30aA/+4CDRhRzir6aVQn+JGuS6Tv7cJrB4lbN8Sc3IKn
ur87aZ5TzUvmMa8E5AUbOc80+bSFwErazISxvLxq6PT8K5abfJVNlmq1pAwAn0H7
CdmVf3y0jcxehZOFH+Cxa1U12DSL8GRAJsy67zoreC5hAbrjTknzhGzutiSpSAcK
Ue78grGZlHEzHMaDrGcFI2ZM/19giQq0n0J58yXWsV9fc+CRJxjEs1ei8dQ5lx2u
GD7/8UUBhIkmP+r/e5fV5mXQ0p/4klYZvaWdeAFHAooUO+YJQDQ6i4pHnzFnWPO0
h0WzWqTTR+YltZxDwoXopNaqMabxhF++h6fvJUuxn6qOXamdyaY4IilZJMr6u0He
QJuxkPhG2t5er4hyBQd/U9IAbwZDswep71uV/jdZPGBDqvt9Ln+1YbJkijCr3+R3
QlYLJeR0aLxlgueH2uHpNuy9IejKKSrPeEEEjlwDuKpFIus/Ge3qaWICjAJklhzC
b/Zyn7B5ZVIN+SHwDLIXdS2Y1NJteASLRdrH9J4t3JoKRFalpLTfHJBeuRxPU+UI
G1AuTp7BK8evAASdnwZ6LvO5Y9NkWV69OP/UTKRg7+JvjJpTpq5Qj+gpS+YBZvLr
SUTyi4nc2Oqw4WeXl09mbAaOvnjtqdYLTKinuQjTup6/J4xYFsuPgwWJ9QCJra4N
CCo/8GnMwdV4opNLOeTfhPTL4hbkmM8ngXgdzgIlzyyGJv75a+YCfoY5r0NEn8TY
Ns8gaXTxz1WYe+cCT5BkncCeRvZhiy6gMoIMQ4Fy41gNKOtjJPmJmsY36BKxOch+
T1elxOXMtoa1kttLrpiWbVEE0SZi8yIdmtMWwROvA6oIfSXm1he9O64ykoBUeKRw
BTIyapr1GbueAb9OTWAwD3VsMX1/vFspCstUp1zxWaAN25oc5GE4M9EH3YX4OTfK
FTRdRQIdClCLyrRlp0TK383SqfbhbfTCiBgiwlvvTzeBxC0UO+t8QVdYnqSVwpFB
M0AI8BphTsyzxsAdKrRn6734Uif30sWuLvC+VYzbahf5HZuPFtIBHsFyqA7LzEGs
HKIAdnf5xK6BVgBfBuulQWLDCkIVajtuJ0jkkc4Ej2DnSYihVuVbZ2nFpIKr0Sja
BXbFvaqYACJcRJJZSVcLZXT0Md0+R6f4wIfCi7l+4HYZsXwQNo/cCepYz+YX/c0S
e27rXTiqpW1nnBvLIpi74JQmKuFhvse8rL3ZKyY2G650I9y9yx5PuTH/zvyd3tYr
1GNiiSAjALcoQ+V9FNQ60/aGydWQ2UQcKQHFmenB+CcUmCl9PM+h7x4+3491u2vQ
ulwpwbYFxWVCmTVvR7xZxUb/fG/VkGUEXtsuF/dJ4pLQMPPqFIGE3QmqcgQ2db6Q
HEXPseywU54uQQr+FzoAikTZYRcTsVBOPDnQub0voQ1YtIYASFF0ed3u6YhJKrfQ
1i7VS6KSH7EdNSsSunAjTAFLw82bMvmn4lSneAKlMWFlNwYNk2ePTzdk/oDjQKfc
aUD+ASanmFBF6A56m4aQI++pf60jEGCdqT2aeQgsjXJY7j7Er6K74RX8DPZKFomT
ULC3cwq7LLG4mpmY+aRDvZGiQV0RkdAYZUS5keej2AIwevW2k/2GAWvAmVNLJ8aB
6K95EUIb+GdhYhQ+SvXf64pMBua9/nddj8RFVZ6KHi7CtzNEBXOaIE+Lh9zjr7/A
HvGHlSarUY4FAo/Nbb3nSUow2Ji/MtD13yNkXxrf7KSbXY5WkvhDhk1JdlO1uc+N
iUxvjb204f+LHMel0uXvMhc81Ca/hcCll84PJcaVk72vHcxvsisevCcZDWx72qnx
JA96ca4ho81eRH0nwyG4GvRch4vYLcandike1mTWwiHD9ACsTfLMZMa7O849a4zI
g+GwvA5Ag3ZHXGM8hobtBTLwoAIwZ+ApwePndj6j6xLDpzYM/pXMvuVRegHkkcYx
WbjMU0bYkiA/odl1RSd6QtMXQxRRn6ZjmGzh6PYRiRsHKXsiotNxXENuEuoiOH1W
ckIfXzv9nSKNnIHcc+VBTWsTVce1E/VDo/vB4p5hdVIapuDuN+KP+57ryBQDJDfi
qPUbf06hMOebEB1qJSCK5puam+fyLbiTo8FpX2ekPR/jhIVstBrpjWk2jNCEPCGN
rcKSMhVg2os6Cb1Wr9sjDJBBTvf6eQ3R30NRvlRWT2ALTgQJJpqtlCgX8U3WlRNs
1enqHnkd9Y69CnB3Kk/NBcLu+Cvc8tZI0GqZSNb6KHAGC4b2JhkIPz97UVfsTKui
WHX8kOXF3a6m7pEwJyIhBY7zqc5pJIEgJRvlYKweuJvgZD25ldQ4jVINMnsrXGqz
kZeIoXxbOoSb1lr+4zct6kNe7UxSVz/177lNIGaaOwT+qS2Ia3Bn+ZazhtNvY9Nr
mQwDPcKTGC1G/C4ESVtWxlkHAJM73SNKIwi1zZY4AuFW5ZHkb5ni9pk42D4nH8QL
j5OXBZzAVk20Q9ELbkgRIl2yli8IchSY8HSseRT8bq2tP4yW4cXU2a7Dt/+ntmn+
ud4H0GPav7iseC+nx9XyET2ruu5sMmQl7xzwI4X5xs7mCWw0Xv0M54gjm/bNnJAQ
secFBusofBic2MuFIv1CxNN2ssYuMIYUOx5odA3tKH1E4O6RA/OVLPPLZVNPWCjW
f6gEWweAWWJtzEaNsMe7aHMtga2NiOhBLdaOJBtADNGLwscRd8/xUcHuPR/QHwmK
jnauh/b/7/iXzWT/uHboP/BV7nPi6gHoLKOyYSSZn8TryNiWXVZRSoGZwMcs+M/0
2uwnthH7451SXt7FfWViZVWP8Itc7cZWTrCXu45U8Z23wUTq+0r7qkGG/fEGqAKH
PDtIAgLYgie4u1Hf9tj4whnln1TEqqLGhPBppUyzrpY9hbgQ9pleg5Ox3csU1lGZ
CJ9w/R6BKFF9dOjnZmc2wuN1Yx+BKv3Ydh9CvWyhnDfmzWKByTxkfMEkiXTQXVz5
Lei+Exf3wXHLgA9kXx74WI2rx1iNNIyxEIg/gDFWxR9olLRDmYSGOlstDw/jgh28
Lkd18h4xn/Bhx3IRI60MDhou4HqbsgeHb/6KMxrIm6BDDlsbAJxUfdxhlYqiznGT
YctueB03CDXijBs8MA7Xca9ehTj3EBAFm7pjF1v+qDkI47xxgfPK5crGrHddkbb+
StJeQc0aD4ZBsAB2zBr6uW5SuTW4jn1GzvIb/y+HgBPZ+7wjTCnHsQl6V9gE3pfz
wGHoryfGznjgahb/AeF2EH8KZGei9F8kKcCTYKUlM2r7eiXSNOZflbNSEwqV4FBq
BxxwXunIYJMryQvWQ19DKY7Hsve8xWSBgBZ0yeB6TcWsB/NAnyyMHmb9N++VwhDB
Mpf3AUHhg2g7yD0hU0pH/cN3LOqQbqyyxTfQFvv++iwYK+8to3DsOPe28rsvWDeC
fF/WQbo6dH/ezkqzvwKiIwvnmCuEd+7qQ00/0zhvUh+H/ZjY+WMbISuMb6VQF3E8
N7eaWhcsxnllkQN79ls7H5FPXR5rEitAZJzc8apx7QsHggdfGTPe30L25xL8z/c6
UMXS1A4Vq2UYPoGJ25S6VLggIp8y4XQ/mtF/o9jiwVl04Y4OI22NbODReRR5Kph6
8xYQmo0NeFWIarooC8+/X4f1rNz20JXjuDudHCFWG0iQZWfLVCHmneP1x//X40sf
KqMmboYbSYnPa0jWKcYCy2qK5b85k2jg4/QoX8XW+57T4/phkVQ252ihR8nFmNYI
uHNYbXYMQZS5Y+niwmU+S+F1kmEazP1bXT6HlXA0yj/GmJwTUsuki6Tz9UXF9eok
2sABONUlM/gV1p/hmiYlTua5Ti9Xb1vX9j01rpT/WszEzVYNZ1+1r6QutHTkjfSh
K4gACbeepLaRtta4SrXg2OvcwfCdNoygNQKyiAAwv2I5hvTjwa2ct/1AUz8ibAqn
znfD9CNURPXyG6OJsCEOib0IpCRAZTDnH2RsFlta3XMhklHjp+rpKvK6fX0VQNUu
fhMo3s+Yef48kF+nfBt1dc4MYT0r9HgoUEtGrEcPO2ZiUW10a79KVxTQ+GxLYZMc
ZeCDPMzdNDlUgTzlSH2cqkPhbzYUpJ64Gv3XRfyeXWk1bAk1RHLYribuSPz9l+Ci
eDnfoUY5o4a1dwwST3kc98m+aDm0X/BMeMfV/R+b52h2wU78fiSQc40QN6KmqTON
V0bx0lPzWLgfcIgJDH+jslXJVplcrnM5GstnEGAqyH+TLICH0Qnb1eiXSEwZbELr
jZwBD/okuFIjBvT0a6khg8Tn0FJM31eGYlKTQK4jBcovG+9u+5sB+oiHmDZIqw2b
Gzza6RfUcI6KGmkWAFm03HuDwacsD5iOocNQtK1VQRPeq2l+128MoKLDWPcpIrfO
f/ZCUSBZUhyYcDAP+6VxXNsaqOdlBbdDDu011/x65OFwZXFKJeA/qpCcW1mtge6N
Fs+hCad7ZwljHYIVCmvcqaLNpnYADOctpKsokD5RCRAcSRn680Fb+boovBgw5pcA
/OEmvIYUE/+7A99ZFc8wivHvCSOh9ZkNrmvgaeHJQPUp6k5zXLjmPmPUVLCRI06q
XqQkYZ0H7KyPkxQyrLRgZgUWwh09BrihHprGB5F2j7MuHbjqG4UIWCn+tZbgB/I/
E8BwcC78mNNVW4esI3fNxcMmiGxHAsIe6cOSrSSkNuijUOU5t0xToUxTrGtLOEZV
dZ9qIA3uArJk3xJAkTGbxdLAr1G8SHZZUEcDmH/q+5bXKgfk7GdnmbaOPi0GPzeF
J4JZsy0YV+kxTm38KAjN3Pr1rPOKSD9JH8toFbGNVo4FcGdbYEpbteUKN3QL8tGt
f/VC08x/kkZ0zeHkYHgpUw23relh2cMi0Tyg3RNbWyRkP5/THKBsXDlWK51X0uYU
2j6mf/1hSVvSC99ThNtaD0u9g45iSFXy5avlY+jaYCA/outtSLCV1fEOmnR09DDP
OUW7N5xQJhzxKOk8yrZ1/e8ebH/w01QOJH2w3T/LBZGFUnmRxNHnM49sjDtOFeU1
PPLiQqpHZIs9CJv+dahaU//t/nMLRvOi+8iKHP3/YP8njDxWZKkaemFpIQpaUED/
Qg6do6dE3slU+D573RQF09GnZJzx0fE7XwLmloCKVLcnneYFB6lOVi79TZnjZEZc
I8U+pewUx3qUhZSQmKCBsPLRcBS8q3F2y24WDdHt02r3ieYGzwfIyFfHCRJ1rSRm
VM5MlIPqXiGSJQtEGuKj5f1WQUkJPCU+/uceRlHFp9ne1tL7V6SY1rq/8TFaH8hv
g1XC9SwO8x0sOtIEKMn+HeJD8oWuJmdHDnTlZDEUkJo4nJc7QfXjOLzvGm8hZBt6
pVTVb9AFyhnLEk/6RUsCZPJidmTTD4vHNAp+EVxX6o4bI+Hhb3QPe+xI5A2zZCkY
C15NIxfysq6TIizq7aCrrd2/NXPPKtDoBr/15h2lg+ncxI13qXi4q2DrAz6ZTW8R
weUHxhXIDDwowtO8YNvLXcMvsXV9B2hv0sxbkS5kq6GXYAtvXBdAXWlD2bB5tjP5
YkM0RnVEyA7LkKit3gK+Xnb0SHXJgjkcDnFJ9Nu5BIlD/+D0MC5Zd3pbk3UXyVGk
5DifEnOBAlHy+wBL+6B8OVqswy4tGct+02hHXShARTTzhnp/2sfMuANbNzyUhus9
zmoZYtwY2oAofjd7m9Kk2XhAcoapbbGeyl1AOwTlDpYSmv2czBHcSobhNVXkTcCL
BZ/Di4z4FMsdSonfqaPDYdOpy/hQdMK+c2X4/DiytM3mpQ4kyvoXO/FZVeClXecf
Dw53GIIdJsQCIv7H1fyLHM4gIn5eHTd2Wo6ZGYA2HXSwkaENiJ3YZ3Mp9TeJ/rD1
Ipyt8XOCkVJ6xQ7z6WvF872CPaxK6s2TEr1cpBAMp9LPAqniE1AUu0qXt1Wi6O9P
NIdvjo18tGme/zs/JvHJmLgoDVVqeJ7GPuoUvkcJZlw1VrSmLlJjDPdBBbcwS8Z+
PlhUB+qzo33lqDB6vGU48R+C1S4lqhejFfutlqraU95HMifX+W+5w6PzNMlxLExk
9OHzUcEgRu+2ootYQmGtCD9LPW/S+U2GdMl71Ih2aHFmiROp6NNbQQXEC/9EKZME
yMI+RSivxgA6/0T45ZYTXQ6qReMCxzvfPsbdECqqiTna7FbfCltVLnGdnb4TCk2g
zYybYvji9pk4EhrDpzjOlznAt/jJ3WwRdE9Sei+KLxxQuIlAa68kiVz+dHWL3Zcw
kyLmEi4gV9rgMUHOPkmUvoMf47cXQ6ayPWF+ztGc+HJmvNDt35v1nfmoCjQ1DrOL
PB6NUDiQvcNitx+lkNvjz4ZTqm3hdiL92TGfkeUB49DiLP0pbm+ULpBo/hQcOEtx
oQjtvp3fI48EBgpm4lht9LMuuGm/3Bpyt9wi3qs7yum4y4BiatBEHs+bkak4GC/J
7C4VMAEczj/UYQV/6SsFCqnYe9zznbG/OGcb23ALX4j2ivRREoydYJS3PMT/gLpx
mc9r8dIIzwA7OKhOmJTb++vOJwFE+oQZO5YC9d9X2KLQKpThVLOVyV3ngSxefMFL
IHrD9t2RzUt+CMWDN7Qg2rbuDxGvn7qzByOJy4aRI9c4VAfx35tmpavRFqMT36C5
OnhLRcvrKmkFy6uXVCKyyqwafEex8eL+9VGBIE4jARx7RkTyBSUv5YdtblueMH1E
9DJoItBOvaMtFbg4wbho8Qe5D0Rbly4zHfWthtbT5bc0GFpI/J1M55upDI40UnYY
qmEwr18cUHOfhcrjV6lDyQQKWqPg1x1pupy2kQSwIPDUvj5po4ppiyeNVOwpzMvX
q7sBr5c739OiuTkLYYNGxncHnIwjD9vg20RO1zYG+siQyt+tLh2Yvn/7SypTaGA4
lXQVUWDOU+gRVlB8swZKDOid1S+OfKkIoj6kRFAvnagXSLt95qOXDMHvNY29QzQp
MsZgVvvnD1dabvYCC1Za7Yq5IJOivAdVrdwXQjffMMbY/GCAG3Z7eie4YFS+Qaa/
O8SWwG3//8rraC7/qYplvVaN5CRMtCANGbnRjrnsm4E7FMoDJrZjEx8gZ8wO4vh4
IV9ge/cwW1sO9iAjsugydsmHMmjhf3MYERv6NqvGKHt/EoJ+ta2W8nC2v9JdyC2o
pIXsgSPS/qZ4zh7/zT5FuuoiAyHg0eLbsVGQ/23zax1NqlJj1q+cSv8LfV7iv0q2
QFnP4lfQcvaKq2TN/l5JPvVpWSiOFVwpZKwzZjU8XnnUDO2gDk82/HUjCmnwk+2P
5HwAf9eSB/OSy4Pur9SplMURWPiETpJY3d5dGduabCFiaWxWQjOgiVGjwQfR4Bxu
pv618d0PIvFxFdYlvgDKAvh8ABiBKwY+cgsHwwwvCbuLB7dcLezlQrv0uxjVuDUI
bmEvw3fbbRCbOzBbJIlAcDkQpn+n3W4K860s18PrtO3KrOc87knWN2qufWwCJD+E
xemavAsO3iWquG9ZoCKFtgzIC2Y8gliG5skg46yxRXVpsinb8ddknwW6HhFtFLK2
SKDwWY4xB3G9eRRLujurmBjudRps6HI70kSjuqlV5v7TB4K3rr8Nz9ai/0jgV+JU
y0gFCU5eTes5dJ2iazo80sDPoZpIkKL9dxXTEwftSiYu6J6oI6Lo5ZRBwq+5UZV1
wu8VD1r1Tv/Z6v2WLjytL+eP2GZLZGpXDFpqstOuFnbRjYUzRTpuE6gNDTz9JkA9
yhC14Dr4vp08PXUaVe9rxB0VhlPwRhqdsO53Mrcu/MqVPuwEiH6/wIs9VMQBUVKe
hmye7708KXDNSxRBkCa7fvg5fvgVd9VVkaAssUrThLSrGQ32CrorMWBDsGi23G2P
ol9nkvGbvMbgfH7SwVUyMEH4yNEQ9XQriAUhbdXvKpBdQIi6udLsYrNgJruCLIsE
j84/RY2DAexQjFu4MLM+rB//I4bge1+xUSKsWSF2GASU9bnF++xIao4BfImNpVmC
aAkl4D5+Bj2axp35WnM+XXLl99sGixGbGh0JBC1Mi4TY/z9MFVUbiW2Ixyyta3kx
N8ZlgoIUJ5lhQDfv9y1LyfrK89G2YkoKH5nc4KgpIddBxdwO/ekmOkQn62LtCVs7
ip+umdc3EbUvxedGqGWrHP5X70RcGqTrDrXE77tvsWwwyHiXyYktab/GvDid2Pqi
oskpQFvhVruDVJe4uTp5lAiHYNpFyVXJrJpCUFxQZGN9sUs3XSQrXA8Lrt8zKjx2
+uX+tWc5ZvwxXdjvUqD8ntZhhMukZuy3ipgdwk/0uzHHH5ZBBDHMZgVOrkdyFTBU
B0zgOtFyTI6pYXhMlxfFA+LeGbyNY8TaFbUKFZ1eGfrTWE5GJ0wTjVSmD9mldiZp
/6Ck599lozjJSMpwcirsZWMRUTLrHl9Qh8OOjZxVzmevgYzhtxwPGwybf4Nj1lIP
h9Su9GW/w8rq6ZPuM+XsY3WUnTEC4X7mxdHkXJfjGouRxburo0s260LG3s4mv9xB
uHCUmQwv4f/k13ZXKCX5hRBWN16hHKYvEuvBHNiLWwkNqnEbHE1TpJjyD8OvyrfW
9PJmyJ2sGjPv1TvUUJ1BeH9zxsR6TnrAKnHmr7MPa1fxY3V6plZJpMgtQsv2FAiY
ikV5U1SNW2N3txu8cp8FkwzMtc88f4b8zGQwr5/EJZfjUam4/2dEZQ1K38fAgZFg
vlsSmRyfKmXjAnat2TFajjXvgUjEr0WUnbTs78mjDbaY66RH4E/RYmlJsBAPMpKW
EMu5ltJpSSZxise6+HhBSlZSTnJcaQh0ZiLE1VJxngJSF8DHDIrzXebNYEwzAAOP
xoenbuQyZk1D1wCwcxrS6bpjYiQyqa+N0M1gVAhJLMfX0WTQfovFjWdGmoD2v2Ei
7dRDlrEH5fDZ7OeurVigTkTCvFoOz/B4HDbGHAf2JCicncwVV8xKM2YxvKUy+/de
aNo4ozVo3xHNpjeRt5m25YQwXnH8C+ZBmOhD9+WhvQ/6IYW0aR0UE4/bA+/b71nh
igkZHvquqY6zqNUIuLpdzBcG9qWYs11rB9whNu714jedfR4Ej3uWgcZ7uAYtvqRs
EzKSwA4HglT5J+M9Uv5041u81Po5B88rhYnLuKwjuH8qw5akxJgW94i2HdHi7noj
HQl93cbGfK2K2TOXwinEIe2HpAhhjQBxTT/WcokgPFl1mnptUaMD7UTV5NGEPhnQ
Mk5AgHgd8JXVaejm3bcHc9GbQPCm+MPzRwKQecnxgkhHHHHRCMV+ZpMgDpt3pHp7
DANASBhvir4qOH/8vdcw1LIizi7RYTokh4ylPLTbU80s2pF6J4f4cfpWf+oupGC7
A4e1E4z5UWDylIVnbX7R47WdaIkZ34B+fvVHBk8L1uRi+KQXUEnIEfIXgJtKgYS0
gGs69YzLIzvVacv32hICTUWIhmztn/OwU2YgcYjxnxbzbXdnGgAWTqFdiSeaO6jA
x7LWpYYCOlpJ2yJfP/c1VEI+VAsnXtnSMFNqftoHdJBX2S2vkiY3g1Ug/YoDGt/y
K9bIq7AdgVBB6S2VgiH/SM+vGC+ZptwNciVLq7FLCMJ40erPBmF1aplnKpDj0DmS
tQcdx1IUsg4oodeEja3Ll1TbeQj04aYKP3xp2zgdWQqrYVTOrKs6Or1qWu5s+i8d
KIJ8D6u8lWM7DWP1sPGgBl2K4qKO+n39mQUz3ZoUDZXLNtrWQO8HqrCQB9EyF7kH
Wg3L+G/1yPB43/xwtNhvDi7Sol09uLJGkuvLB+nOXC1HcIw4ICakRJO4tz4xHbOp
+wG/B5eISfWmswzDFmYBfgCmpxA7ZOP8D0S1/183g7CYKsJaZ1jy/I0JNCykBMnx
ScqKlwIunA/mqC1RFgJuQAHj06j3QBO3O/rysbbYOzoONCGLdiGSQMzY/keBCPNL
oECpifJnBGdloxdlCo0KWyR1INIp42eeE2JGtl4eAl+djdp350PkM66BL8tX4owt
9s1xZEGwUVyCem8OT2SFlUXuzRii66kVUhH4sKVuqLEPEO0lCJlEz3eJQPBRIMnC
MXiIDl/+QD6YhQYlf1vHMkKYUWnn8kxy4cys9tTOeMTO6Py+0N3W9sIkYJclvfF6
E9hBUjKQijdPwDG83Xawq1SIOXcB5D7koOXWSK3RbPUDXSwm886w/DprPi+331l0
M47D9oa+XI3iosz1oGaryNTuM3LwqEgO/5rQUasvhVHD1WXH1rOM90xrqQ80eadl
2UQR6reRAMwlLNR2/NSSw7/4LnFxFe+C0o9MFZUvILFk4FhG2XdZJYf986YfFksZ
dAuZDKmOZvIXowNYBhuB2mii7cVKazV6xut6NStA6+huMNAuRHWWo+YcVVWfIP9w
0J5DnroUdsq9ewUt+/XaKruFQRfmqc7twq/eO5f4B52a7u4A7ncR4HRV9PCwuh2V
V7y/LkiiKGsmu70hsGse7J2Ci88/yXLjUjed8tFstND9YVcbDhxiniNuCCUrP94k
TxitFRXUOVpQtMaJZE+8QHFbAKdSScXTtr9LWjTrc5TiecKJfma5NTpt5///LXNJ
9dA3GLLEZSyouWMBsKETxIj+0fTRh9ZgDLhKcRFeX3CoBRQr+IiEEzk6M/eckOZH
ltSybVTUOiB+W2flgcRWpnYd7+UouhPQqaBu1km43FT5SXhvkXVRdvodH73I8XGH
adVOIn8lmozSHZcNCHdjR4sv7dPguVmZpYOVhDe9OYIIWuyVb6+3wJ57crDjbylb
w/pGgySmbh6jtE46Ur2/4xhJDMg9tAJ7hgcjcm2LiGXw9Lyl29Wusj1ZDzB9kIJq
SEmKydHdX42Mgzme5/Uq0/4ScGrCNzAqf0cXPqDQ8DUpVh+FZJQJGcALli3rUVL5
Hy6ihm31H/TLwN+C8dAQb47NHmE9DEHoWTp466GVDRpHhm+ciRLPRWjFO4PQ4yld
wPM4ZR5XMXfUzj2YWyOYlPmChi3y42WVjcuob9ndBKUqSvTh9opJ520A3YaIwuHD
vV+z+MXF7jOiQCd5rX+gJVIpq5oh8IVf+FyMRPe3A072xgAkWHfqJM7jnBAhSuov
rm+pIMcztp2qigHE8hQuZ76I0p1ubpn3WP6Wz1WYSLXpR2OVrDKUAEZoxXXV4RVA
S2E/qrMAIETH+rmQGA3o62aJIsyXB8ne/V6jkh8D/k6pwzlozP19vFsCrr9EdodD
N8M1Rl8OD4Qv2xsH3VibIIa74FWjEc93RXNLOYFOGLioVEAY8SvIn4KbNHeEYIdz
dTC+ZZ2PoKfAyfH1baI2XJqW7TB0VmdbLnmVrqgBNl8FwyUAzbE8tpp8U7J7wjKi
JyqlMCaO9f35IM7oj9VukHmLB81ThvIutPYjqGQSI77zUvJJWJgGOm5buUCJL1cy
/XLi6l7nXky1AY2epBtFl2wXRRWvl63AyO9sEpGOuu/gWcnhr2TE1GvrzzpXnVMs
6ZDHtxrRbMsjfe4Stj9fNpA72fRbcj6dZx8avYTuulctxfsobvZ5VMS+ibIMhShi
I42m4tRPVljd2OKGJfBTR0BsY/ROi1FYV8qoiSFYiEcT2GXoGB28VQGKg3pOjlpT
zPOD0P451pMz2QkrBodsonYceHejn+fYLgjfzp+HzDaX0mCczuiA0dvYhUyfaXuc
UB0iX2ILS1CIOEwzz3fHjjarSGxHB99iUvTcLh/9OGvW53nqygvH9JpeSU71ccve
RCsFTrZngWjAJWF+XPsQjuXheMVl+FwMCagTrvS/7uBPr5gm5bI/Xt0lzS8NstCt
mFRodzzQiKcXa9oyvWOSD1v84ux2cucAy8i3H0uGVP5m4nc+12vAvpLOW88ykOvB
q1ALlo8eaEqJ5TlvBIe8T5YRDhYMucZg8ozPRaByKc006IslA9bjWW10TQs9NCDR
Sxp36jgFWSLqPZWx8Mi+OTx2GcejNEkDoKE6fzSEl/XmeakjunuFM4SWYkRYq6be
i+7bCK7SkoXyGHrPHJ9h+lsfUJpYpaxG8w6MLqZdT3jqXi6gcJagwz5UGcj8kXvm
9E3dflaS5GmvgNXjpu36HbMer3L8uLhpjrk2GqiR2FumYYoZbIaqnRTOuCjgdpMj
taZwPkCq4nHcwcW8BH7bn6pVakf8yRIHTa/Mc1l/sug/pH8+Nn47bRtjXLYTb3Tz
qW96aFub0i95itJsQv/N8unDFWgRI/jYHt5RmFtaJX9zoNYbgcsXcrb5C/R6XRp8
C8gRJaPKRPtUYz+cL31bRe0jfwmAcLXV7BsjLvBjdnaabxbEIDKhHYx9Nx/WEY8k
81TPQ4Jp/v5kqTLUoW6z/8nJvsL/vPBhTVvmhHXjS3uk/sSMPN6XMs8kdwdb1M76
0uBovC0U31h56ZWAhXF8jlN5vKlrqOI67iS4xVSzjceg5+uufx/h8Hnp3dn1Id6S
3m+WJQMdcELwrW9mE9DcrRAbGsoIMuDvhDUbJiYEcRrQFiRNNMWAJJVjioETydMX
w+HPIvmzzgwtjGaRYSRkOgWRf114B3yD6J+32d2sO2WhdifmIWPT6Z4XdW9t++HE
Mz2RsqosSfNbluwet/Rr+9Tz22Vp+4A55v1a7Si4vymJave8vtxTJtglEF95MdGi
HrVNuMU1gAwyvpI2S7KVRs8tVyO7aMjh9bzUMpovh45PbT2fEO9zjvtkhcRhAV4X
q5lEv9Y3WuAFrpy3+w+ioONruuJoLr/Jc4wGH4Lm3mFxadOYQScH50F3MT63FkDh
rqzglmT5cP5LxHoYStm3qWl96UZf0Xdz+Mo1OWFcLq5WWJRKAgim20j1VPFvsKXh
Z/tEEnbrFi5C0gKpmsh4nsALUquw6rQJDeBhiRBjkQRuBQyGCBbEBAy2qPcw9YFt
O3C3MvDa+Usro6hU48CWUuTUQG+Ukk6DdwT39QpJuBbRgKGpjjDCOCR64lqKjkF7
WKP8tOobMJqduHsMQB3W3advsnctNOvC8PiheJNba0l1eZqckY64YcGTS8BC3RWB
pmWZps9kjGMY7Pa9UxSFEmO8aBSNwZBi8w6iRKSHYL+z9kgv+sh1SKK1dxfUQ/dJ
IZNBaV25Tds9Agn05ql6+WfDsgR9rXk6oV5oknoYsNQbHXMmloZDqPqR7SumXecg
6rffd/ihLCW3ICliWNtuqJcermBDf1DrMyZvxv50BGKF32d7XVgmvTFU2ePuog36
z/mG/kLNwXFHrAX0PSU+a8ndIpJz3zmt20QU3iqIIBqCokgZmBGmPYOnDg/v244A
rQQADOuTLrDZ2ZHqvvtPGzhQ7uMWzqdITgvouSM9yP98ya35Ew567IEONI48yBH0
akgs4W4SL8FnBpwVkjhX09TxzRk6z7AMTFg0XOduU3mWzUHDkiXfb5ymnH1rqdFr
GxoIfO7s4rM/GJLa1OWiJOnmLgevD3pU7Vo4AK3ffq/MmzbAN2kwOXk32kqOIDKY
Gzd0vL8obyf0WhtwxX5PGp5TjI3YgT2pvsoG4MVqEb22z2/Fwi/U6TYnzlnemjgq
2buMGMGzBV1sJq1QiXfDzAoxqRHeJUUm1198ngRAjmSTl6vLHX1L8RhI+l/cPTZM
OLaWbYfZkfFxyCllQ5hbl4xD7ILIVk5QhFXzdIy4miIKSsp4PKwHJWPTMARHy9ZA
islyNqHhjqWlVR++P5AW0gHuLUA4PuCBqEMtUkO+HAqwGDDMQdTiTl/GQ+A2E4l9
aYzextcUzxk4hEUg4RolpETfNKnLHyiUSS0oEIsJ9b1CfmOXhTxRfLIktao8Gd8k
SDLzwZe2dkPSZz/0JiPvqlIAFKBScqTWJTCAK2M6WzELHG8GSI0YdmZYVmtvM/Zm
V/lC9OXV0OwhqiIacktJanz2iQ9Bg0f0p4oEv3t9L/sY48ABTM5fbb2KP9VALOBV
t/SURlr80eLccZSXk8Ln7hE76bKcUi2M+1IUMHKWp9X39ZiwR1cfB2mW5OqbGJTa
77LSGRnvuFBvmHrBrF+WQx68KXcq8mpws+lXbcXmRSPaaTqRwHL9goHaKY3g/GfM
3JWuj0/dhByktLzd3DH26rPcgANqaboGxAxGop/xU5pYNLD8Z9GSzXbzYt8vj21X
hiY6/ZiteEUUyXDuzUPyrFnwPdukp+JH98WeN/KVL4tIOlsBhGEserkoD7bKl2Xk
YFjoGmfFesTOE4avI8fYETh924bm963kBsZZWQNa11OFcie3SMom2NMWQe1CYgWK
tqnaGmxxhUsscDNGE6YecxX5Qj6D4XHAqCwp/ycc9CfVCBALjcjfFHF9qJpeCZ9e
wV/aAT2wUq89r9L4NcdUj+mrnVj2Y+B+2gB+Y+jQhDRwDvvj3GFBrKUZLqh4MqUR
mGH5zQhllp7RuQVgTe7zUmo55o7X05/+UFBKYQFqVN0S783d1XKEe/em4shCgoWz
xFTZBcLlnrbPlYy58l5RT5xz8MP4qpZk3RToHF6fCw7RSq7u9f4VImrsCF7e69WI
JqXAmpbNLPT8ykFmlViDB4MH7zCM/awUTIJ7gn74t5vFL5qiu+Fbv9hCmwX/EhLF
YgKNpiXpRvdlSx3L9HKZ6rnGjTZgtO6aWrMRsPgBsGA3cvnT6EOYlFZlAAMyF+zt
ZZbivYqiGa/0Nva5dWRNQMCYJ2h4JbJOs1vN5C5CamgFyBfLHWHaLg0zuLpo74v6
WgggwpG7HKhAiR7pJnX56WmuUGGAgr3XG6uOU8Z/qCuOImw/WY8eMrCAi5tevuEI
abZmaUjWgLI3VKOkEAlduQ0mWh/KQzCDffJ+g7G0pdto8vgf17L+iBZaXqoUEOcs
1tTBzMLJRJN87mQ7QG7OLFNsg3hCjrrZIgX26omxkXYWasR0IPoBc3DhIXeKaZrF
ZVDEp5zbSHujskJFnqTbeHtrd9dxuybIfIi2q2hXlTxHXL3KFmyrs7c7c4yyWi0Z
2xwiuwWIdsJP2nqS9OTa7HP8ALaGywqK+uFmaPsMFJKD/3DvWyVTFHDzY/Hp3s3F
yfDUdWr/8ttGHHqYyMj1zEOYancQS77MU2ATEwTF3JIZcBMoSO6KPMb3x0WWS33M
TAx4ANO0dyz5e8j2shbEbwWdstWRmphk8WdiwUJh6yONLtSnZpFbvOACxGvUawi3
o1QCTktXj4uz5mDGqRMeOhsj4i0zsm8UGS2zSovJUww7A6XNCuEsf26VnhVaPASw
Gr0PI66Xz74hcd10HIrpSlA3s/pkqwGaW5ArBIe5CAOZdm6+t80z6gK+2Aj7QQVz
o6yrsUDbqvrso3JtFj0QDrOOWNauRJuDu23yI9VLqBEkHzFwcMrjLhpRi7wRQIDJ
f1F19x+b6JLvi2ZuOutt4NNjgGpH8YQilB1IEuhDHXJsugI4y0TfjNPaqJ3DgQP3
MQa/vWO2g0nIGdpW6xctuPwfKgjG3TjYMfU5DysAcc2nKdloAd4NiGoW3M4K4/gY
6CxOugeIymXpD+qFPwTFrkRn/Jv53kMGM0H25lh3HsWAWN/Nnb7oRL6Wi/mPLVoY
tO1UzsgPVZ7kcOWEQc6ih4ilLgrG5LeP61D4HbjCAaDngfy2Hfgers2+LegbPhTF
Mq53O5Mm5ZmDBsLFBVrDOAnXcZLFrAsr2K8xshDRTgrF85ApnykbOyk/9YepypnM
fbjzy6L2TjzGQHLHl4br2OVY/EiCg0AVV+8JyI/H/Ahgd7PfnWZYywnKXphjMu9F
l32roEorUb2nVgsf3H+ExELUrWX+BTuJQL0eKkASKtKfdjqFT6hHgmT5r0f74UNU
UYwDaRMfz1CxfJKvIeNKzR87Y2KoLzCI4gP2HN1e4KEypVP4LHof92AxyoFT8lHk
+ME4NO+WUNAcrSq97l2soEOu9qlZBgCivrW4cEUH7W+c06RvaewvbzyO0ntB/3A2
LL3dEfGWofNATmLnBxqpl6cIGdJJLP/pyoxES5B3sYv2g5taes0SLFwa9c68wr2A
QCqjR/i+CnHkGbkpaMzLEShQb1ab7uUKyYUVWe0Yp2ouUOPDfMdQ7CRsgc47Ew0e
/JK9fCGSTymmlw05twlWsUxhg4Dxe8HCyLKepf+nG2MOL2xzX/TPGjB+htnDgU1W
aMoD3KZzHzvQh+UUHLHCoW8Zg8VCiWNEDj0O/mGZRqgFy6VuCNmgiOUN0CCEz1Pl
YGhqhOV0dCyQjeZJUOC3OI0TV2j79MPF9uU8vLPQb1EjChYWkt/D4Z7n3ygMcrLR
eEfwxXhWQAsDZWII6ub4kBPohEne+3kXuI+cWCD9sHQdUmV9EDCS3Jd11Pvc4Z3w
O6mj6Yz7e0XJBn5BZTtl50TwpvHLpXVj7MXqdteJu9MkG2tUvhTHiPhh5fPWJQOM
lY5tiDuIcNmCgbOoCsSVxF9DQb0JT8HdFXvn2bNCPK5iJcdCJc811IqtGJhd5RfF
KLw8wzrk9bb/ZOy/evXAO1iKESLA5fA+r8V9x2le8qN4JqmTS/hWW9taSkPjjwgW
oDKVN+fjAoTgTdxOdj5auw5LDh9eLTFFlloMlvZEPTEUuuz+lmvNC4Iahk9kI13X
rnI687FFEZQXGsQqXtELfcQoN8cRgZOSkcLy5jiRsPbwJsDPwWpnmPOr3jH5xY5a
HNK7/2QeTEPr4vXFkt9keQod6/bIkyV39PnkgHB3QiD28biMC0R9d6BDXrjmufBJ
D8Y4gQW7ZGR5XVXdjVky1k5Fje5xGUgCue5ckF3jT8w/RmX0/FgM4BbaiX9zygmu
j1i3bTAr8MdeyGjQ7He17xdbb8YhsCXOtdMUrkDJW5UxXEkJ2X8ZfCAUhJbhD92r
WKJqwy4LSyz8cALtTuAFGbO9Dq9z16knffFu8qGgVDKGzDI/bGvampCGeEpNdF8Y
hIF2YZiEmOk7F5jZrRgaJdxNYu4b2GJznLMgmrmDRRQOFzX42bOHcaj3tBYtdGjb
LiHOIvzSYRuTTtidWGJl+GlQr7INtomoMwFDT8+dVBYViorwmVpu6cokOF1UdNid
/b7X1Bop/3Z/NYCePpB5J+r6t/BAU+Xiz9VH9yopWSmpLjGqkF5jYit1usEVMFl6
oIwOZu9JUoFmTUL8Ztk8PkVrG/u3+91ryIJdCDZfSesYHf4lGZbHmRJVtEUzwp8c
yW8JIKVLgBF19CBIIzfdwGB01JF1mKfKmJUgKVAOVzJ7v19Hg9EKp38T2Dyjzcqy
e54iBqGCbb55vaKrrmqguNOfGl0f4e5SrLe7hkSE8Q5sKvjaEhWLQcMYdN/eMav9
xA+KV158Ke7iAT5XlBNG/VZ99VRqMkkbdgVE06HQ30osmy2NyJo7dq6xnP9ShZNz
Q53gh7YD1Bxkr3VzsJdM/Xn22fVrygpq3p/nqEHe1B1Zz8tUM6aM9YlZD2/epls6
fYgCVZgTFFPDRZrgs/lQ1b/LwT0N44IENXyS33791rsfjwSjmoxyyIw5Lcs5ZT9j
XdrL/zn0ajhSiSv9KO6KuV7xhcVGe/Amp6MZALtE6XvBb+vnLgfWj7o4GUSowqgs
vMmyKWeOvtk7POyXic5My1nkdaIbuvSewNr8sOXS3Iq7TApKEEDyD7XkS/3YVuTF
+P1QqWw9FwkRSv6kXs11AhhhyAQdagpNYzZGnnDNR32xz8GU0gg8MXFtoYyq0GOL
BEUDZ0DNzBcZ+z3ALfFivvsiQg+asc4VWgIsVELhDiJAwuSnhLhI5XZczMP0XFRL
PKGlrFZ1EVMm+uyJli8pq8FWZOqulWIQenn8yvSa6iCBYxHWMnmiMao/lJG2aVBf
t/i4ngef8G3J+UrknJ2HIc2JLffA5zQlaJyWRvT0kTHSXQczbFqZPexMocAf1Yl5
jO5r06NVgDJjbFaLSyV+388ux05l1EtnXTJqjPwIWPFdwmzJleH909mrx4NrF9Bh
Hn3by152FjCbpNTH55JPkIG1LU7xGFuawnVwo4nGBDgJNYX9njeGZ9zXZ6c5KH6W
L0BkxCe+UJaPR0011fsBRwXHex501xWPLIgXdWZXlwbVnDkRGe48reX3MVufw2xF
WCsRljVvebP8ZhGBHpsRH6kv7VQP5dfp7B/ggMR45BvaTGsCRvfkQYdZJRtEKFdw
o6OwFKwxq5ZSIOFlyMmls/lNVE6xTPdH0ftVKghu4R8eE7Odg0vrY8JPBOcbqa8q
ghJ7Q8yeJ+sATaSiBbuNT0zu007L7t4CK+YgsnGeA5Q3KcVpAginiFE8dR2c9xvA
McrRrmi87vzsvo9UJysxfeP/JTnrZcXQZG0wUeMaAK0yMLYBfINJBsoG/vsOoGxv
4ZgiOVUh8WT5qq0UR4+NCqmA77sa0vWpOo9oNfW7vchI58Zs+YQwEnJiAbc6ciXp
pbFYLFJWrkg5MaHEEgPyRTgR7TA2SRZTUBzWNYoAqSXIQHW7jPJ2ZPDluFJ20B7K
7CQcEze1Brn66dtI6HMOuRfRr2vNWy4AQJOecw5iIA25uUokZ+S9WupjMYgG7KxL
FKG/dcI63K5ARm0pkUfAcWMwVrC9YGPBMm1OpyXGj7AAweXSeC4TnrlaNmbYXMDk
ofjLcNrZZi7LqFTGH3EjP6t5jN7Q7rLckEUoXV6fWdINeQ+smE8yxlJc1z4qGNzc
SIfqii6KPuagPQhUCiaoZlSWNl0uEALsZies7EP0aQCO97oacjQVNSvOsaDGF4Er
vuhYdcKzTvptw7Aji9g7ZN++B1EqbSDlT1rp7qGrBawihBxzc84VjQxZ8K0gKQ0R
jKbG0vS0D/1zlZlMUSQbwTfVnrKA929+hfIpIs7si8xDq27RmGhfTZqjOzrfo/r9
O5yqZ2hpbGQ+1Fy91dexONag57aaeR1Dw2rZYTyBQxm2z8k8ReVIyvEx7W2zJGsf
3ZufueJQTGq9P//mgbUSiPSbqpN/vs82SAW4Huu7i8Uyg9Ctju61WOlnMjNsKokp
WG7g848F5pMk7Ax8/B4JokQul4IhheS6/qll4otRPbNqYVpAsM4n98+TXIf+SLQU
RjjpXJnK5coX0dnGmXUSYWK438fRfJvHmJGpvvycIGBqjJRIxjuXe1fMzL3S1Zzq
IZZJEQuiqoMZzPN4KKDgX/P7M21PMdINbOUyeH8e66FTw/ZWV1dUraUUQc273w+3
ZwgMG0PwzIEafHop+vgKCFQkJ+leBNJTCL6nXXmTpJ0pY70J2QxFKZ/XTcujhg0g
Me8A77P4xfjCleumSkFcG5Q+VShbXloLkyEKezzautn71NzDelUHF9cdc4ikBDOc
6oYijFN6Z3/YzGhHPw4w0yuQnoPX2QNopMHtan4y4pbhuq1yNWtSIUCL66OeklPp
s70kIH3xgjHXbmaK0QrBIc1+6kSyeeduxZj4IFZYRx/M0LAbcn8WRKS7Pn9MUX1Y
5WlqU65k1VcWT5lpWpHsZ0hFA2mcPgwEn2u9lcg0OuewlxX6UfIDf+Tp0EGzbFLK
BNaFVhwFt/+Le6ZzuimNg3dauNdtfsp8e65Oqb5cmrQu09vmDMxCH4O0xIoMJVRn
axlrbJRaQ8+bNNn+kqPdTJ9as8HTJOTl2ETuvz1C7W+fNvrGPvIU+ykPrE3Msbkm
KKaYEhIal2G7F7wUr1UnA1tsRK02pPr0cUJ+kY/i075OuuC9Ta8+y/rRXo7oK4Qz
VgZRPjn6pYCl45P+tBap2206juYAL6iTI/w4xR0OLKEMnw3WZqzu3lSe4sKIdXwm
7ECYMcFBWdGI3GhdAT+fFhOFWwYjdoyo5M3IhJdMcmLd49f7eDZEocaxQXdqOiuy
O5Hu1nkjde2u2Qi11MvA35WHg+2gJmgPvKeGa75wNQfkmzZRX+8c/MHGVnW9AlAk
scWBXfQ7N7wcgfFCgP53GTQjdcsFX67LwU0qsYSCovDqtKSZPAJw0meimNPTYQ+m
R7/1bsZc5tS8zNeIZocZ0DH4AlcQLks8wD3hMwiEOX0KWRBACKu0gb7KgiQiiqOB
LpHyPCvXSr0DZTg94uJzBtLcdnDCTPWPrdoB2kBkOahm2ggboT3k632K/uG4Cqct
sERVLyZt4/fAptyqkXdfuIHhQEMQbpqzo6yrkE08Cj6xdWnpPs0m+C9SvtSQrKoL
bHbu8yv7IvruVeUUb7yT50c6ohufwVnASO7V51m+1l8JQRtkU9EzjN+dRdKkwQOz
UdZYrXP0/qWXXJcnGqQqw9/BwhIZdoSSsWWRQ92lw4R14BwjF/IYUzW83HEh4Ek+
cBNjbGdyvA52mVz3MEZX3KiEOZiAbJP/Qn8nhIzJlqpQQRP2Who4Bq/WMIsSn6PR
cwlGGa4BNjUr+AyDgM3CW5XMXPkyfp7tzlcZ+PXbGyFRKVKLBvC02H/8wYnGNOrw
HIzuFHMy4MfUSfLvmU6R4o+AVaedYO4s/rSXOD9OV83pGtqCMe1xLReepAZEGWwN
/iMcggIcuhmuGiro46VevOKziWTvcuKiAhm3eDnRkS8kvW8Ij/oupbh6m0TUNeGN
wY4peHOukvCH1YFrAmTJ+DDjoSytxywSeVfb8+AX06L+lvkQvuzgKBQA85r/tWOw
B3Di7571zHlCstSg1LcTf+CQA4Zysy8DdVkmVRfAk/j70kDZN9f1Zo7P6tFdEaZa
sAJf4MbOG77u2OAb3IwYoKBlL7dTwy3dzUwMx4uj0wM2RN+GCTGzvW5L0kY7Ri7m
U42Hoh/rQUEZwRxMzt20At1oFx6s4xwoK1yVOG7JTl0UxbU8/TFhj0HKmkhWnoJn
KiIHq6mliTGeN0ojNGHEmzk/UqcTMhhkDVkuGlP9tIC0IGpA+DhGHuocQvdCOBtu
Bkkp6zKyLMIc/xwv459IaZsy7NNOb9qzO5bo7zXIKXh8ooM7N7tXJhhf3cOulqBy
a6vYBuShxhCCDDLWvzHqWhHA1US+sh3541AmoNgmXGLktj0ZkNJj+2ALmTuPWhzH
/NIFh/D5SDWAHtBpkz44/xgl48JKiPRfEgvfWY9QvFFjHXAWOQ/ilOlpqt/7Cjf6
xHuSc8Fb5hSIJzBCgKBIz54GCfRTELznwjxsrmX9XM3yaU8yQl2z9d5i0ZuNNujY
NfMt7/VsUyzlM3YyQvhG4b23jpzw+fS8gAo5K6ZeRpWdauhUXbvvD9tu367USsvy
+jxZTgVxBsvsKnnL7yyXa2mPSoyVwT/hveVl8uPG+W69WWttlZdKF97ysmOW2wp6
ThuA3Bp3KN1/MQ+IEmCHxMxOG0bU6MBLwe6udxmR+RJKpiH/kME1WHbJTd9GHjoO
ucjstWicpy4Wvhw5LU8NrtVGlbVfpbCdoOSzah+yU1DBiuSqUfJ57R1xj8oSHYMk
DZHg/gaj4J7Uw8AJZTyTJm+1+J4i5VMNy4mJxcnHLXPV8O6clteziJy8E56MqTyT
i5RokUschVLv7tZ9S7QfobU7krftZO2ns2ScW9OFyFsJvDfnUtBNklnH9I224M9R
bPlF8NRSLNqZAndu89Njb52n/ovB0fE8juG9IJMT5+T9VSFBoFKzalbaTWIjJJkF
QDW596gslBhX79veujKT/MD5UAm7ErKf2TdV25HUH5+C072ENi7FQUsFxWoZoPDY
AGY90F+Fq/UF+S0UXuCv+egvUvHLxkLwL7wOHrkB8hayyNz/rpVuX2MXQdGt/QYs
18oqEOZh1rYz4NNBXvEjdg2hyuZ1K62i8ulyeAxsmDMQ9s0JqhQdYX+RK4lvEK9T
NMzaEWMzjfebSKnZm69Lc/APvEkcJNKDxSPDOK2cHx7aGhzKPmHOOJZbta+zOwDy
PiKk51CLpE1Tj420sWzMsgUe9fhPCJpfkAxAc1zMN4D5Cqi1BMHnqT7it9DNqYSR
7WsG9YPhPqiFVijH2R59xG69HugO93nSqyG4mkVzddL+XV8Dbj1MVC3jf19xzAIA
Uc9PjyNxzMFP+jtU2xLPA4wip2r5JrbpH8VWfLM+1D88xMZj9wjkro1DxlOl5zSG
akA/5N3Y/oBwJZrQsH8XTmKUTYIXOE4McAaCcWo2fOs3KMPPUZH068q3CZYIGaBq
np8tVCD9W/H83YQhqBXGKknj+PxJvvhmtYdybv3A2Gqm8hhJTRyFE+JKFSnrV6nK
hwO+sNv+P8SO6PA6nbvZyYoxTd+aaLNedRaVGthLlMJXkT1DFlbgj4VhHohCO6NF
hz8tGzqktjcRh4FOz3TOid/Izkm7D3pNwac65mnPltsA2TsgMhM2ATUBLW906xiO
OQ3x3PwTuXL1tPZJWN0LVHDJOztkMDbCc7q97raLYK1vGEuB/LkaWiBwtp+C9DjO
WYZGsThsw+xHBm/vg5Y3ud0yc86/BwTpT+TKwHKchhAf16FeSGe51B85IhyihOmO
5CQl5TuPuxJJ4cxOW7HKwbhAIvODOo1J62amLXKHsxLOQqq1nhX88qatWbEuF2Fs
kqWcvptRdALBXAUvEZnYLn0LyvXp+fogWcjCecUYkhFIQ0Mpb+uUSu43HaPkpKOe
NMSXPSwZjJycbRvZK1pB/4xxjFwdDmmzLQlNJuL+dkGCxfjSCSaya8DQLaoSy9Uc
4Ej65ZdL9BdwVF1I8AVkwGZqA3aOa0DNCZakVYRwwYXqPphFjrDDvZ7vtBpwB+VZ
jjwfGoQt0AiECN9tXBYiAMOVEYwPsi6V894vclZ4ZFYDA37/P/D+4Scij67EkMjR
Kc/XxJAmHRWY5Ex/aFbbS6X+a9UoC4K7221jJIXt80V55AMofXpUzoY28Z4M2UkS
vQhVNQXlkpqb+gkuvijZs2OvrXHW0J9+yTAYQseIncJ6vEF16QtvnctAIK1/UeHT
H6y7+5eDE1Is5g+DKKYRofQ6JPyLCQiRTENiSsDWlmw9OCpYKTuTT2xYA3FYOC/o
re4EBBWXYy9UL9j93caBnzhbe8CITWERZptdZF3i/q+44V7OossG8TUXZ6kkf7Ne
JrByUztwDqDbCPfPgTtVjCIUWxt29nPifEpR+VYoY/qAebNUkjmojjqmZfoFi3S5
DnPCVICkb8acvMsovUxAubC549ac3cx/eZ1CV+mG5hP42hQUHei9mP6imkE8fbJa
eife54WZ1oD1hFzMugNaakxgw3YoZ4IM7n/KBnbSEZx7/1A5GC2p8oH8rWcGAtH3
gnhSzPsDCTLVFglAAvvMFy84Eat4Xo2D6TB9g5m5bh3+88LgZqAB8sytbIDYI14E
lD7e38jf8uBULCcPn1mKV8VXWx0A0T79xRyBSn/2P4nsodjO5mHXxrQYIdBPqyCW
QjHsgH0GdSlPCiE5lJWiEZSJ+xpYHnPkb1mP1XjvCfaUI/Ok0UJPhnh1i1tMOh+p
uczetPYUbNLF1A5y6bwJtNVzAcrMwEhh4SHM0xik5wr0IvA0oC30haHpaC1Udnbs
PpdvmSFTByd8FV0Z6jmVrEO9bsYkR8KtAochZ+Pxz/xHNhNW7XQw+M8v6g4hfvJ9
H6U/5WH163RuAW2t6GNo7z5sRPZolM4bXsH+3BQYCXLQEXV7efByqVOc7BNdJ9pW
1TH+vhrwRvUGVCfSUbQ8wAIZwdjaY6uNExr5EOSAFP2jkNCnMwIvSC1yJOZkkD5k
W/yWL7MRjNDFsxT/onjD+Q91TjTV4NRCZmPEM7BgTrhJyHtvL+QSTMZR2ieTh+Tg
nFcVMN6i8hEyskum/W3cwYDtlPbfm8kajMt5J5QWukipXTRFvfR5g01jXCM5/L5L
VmisyJy5Vl+QnyuyJi56fj6FUQ0GTUEiZErUEOg0diOGY4uDjA25TGtH6/OTwMWc
UJUpyGykK85w5ALcpA4SWfcJDeKlSkAtSu6f/kYe9odBKsN6sj2YPuxNKoK9YIGB
dTPWNxxWL3ksrBZWdr9TZr2Q0EVSgGlv9nFyBW2a+wp5cTyvONiLIlFyQdGhFjwv
LOr5eVSFC4s4yCecykR6D1VtH0ize6ecNb+aG75/fUB8VmQRVovULQrFt3olKVo6
O4CTzvUz0AQS4gSVAPXM3MsTe00ytLiPKC13OGdtpjTqEmEKHXpFwTdCsEDK/6R7
GLbmMF9jajEF9JfWbfKrsgl8Imr+1R3Sng6ZE4g6AldUTA6RxqBtT/uv1J4mT4mH
b6Fj+WwFcbFN/wT/1+HE4JSUX2bW3D9G//D2eHkTn7Px1vrrMZRwGCNzZXfcCQyx
v4e3W4jQ8eA0b8CrgsZu5Wfgz7B6qXsA93CZ/8vayWEUfwxVfhq1k7LDD+PAVh+g
iN0HRk1YfPeuiYDoT2nJBDBmzYS7odJRveemtLwOIHUYt0PmU2NdkI4oHYDkBTIP
sLI8JIkI/ZIH038gDmGokTJyqn+chR3VXw6cwTF31Z9UPWSJK0dJEQZjbnnSo1eU
QXz8DaC+dXVBcEJ78mWDv6HQDvX+78pzyUGMa3jICDaDNx3v7ruC6WQMoYHsui56
zkUHBm4+gmqA2XysKrlfPuZ2Yh8TKVpvm/u03ixyOOph1qhHDyvXPeG1SAAG8ydG
s+m0JRrQ5ej4bHEJ0y6Ag8iNlhGgPoj/J4ODqBkJ6EulJRsrWTRhSyUNug+6jGl6
Me9uGUR0TaQPhXzdYXje7UB7nLId98NTSHeyCL8Y5TyVDXTQ/JKc+R8Ur5xJKZly
P3MspPfCIeVw3QQxW2FS6yys305haE8Ve7r7U8GqclC06g1YPXRfvJOa1zhCqJe+
sDuyp4cTjdBkW2rUY6nreAgT3xABITayZY0RcdV7UC8J5TknEgGTZfXxUySizRWy
b3BFRuON5Z1f82z5QmBUi1dKszpg6DpDOB1FF6+RsKT4Qht6bmevkmSuRLYtGxdj
vCCaNs9mG4q7NIWV1Ac9oOE6Jw2lbgWC6LjOtWjjnmNmF3JlfPGFCcw16mvq7D5h
Wc4rDsnpM5wTqGFY2xOsBMt4edImN7ZXrIvIBn1gCj7YRU3EuaXnt4k2EvZbKlS0
9dwlFonoSUU44rr4gmQ2eirILRXVsiXUzQdwTTpD7cohf6rPR0LXRrp+H900oayU
TNRZHEcLlTYh6rywzogdNbZyFyVhssi1KyQioeXJV67z5gqsKe3YgzKQC8GWphrG
IT4HEDmVayb4NbHUqj3SGc8SfHgeU0Vr669vxgOygUgcUIfgQ5PoxcQioSkoOJwr
ngAXnonwH+zHIGsTAn6c9p1/8objRGz0yHoYaU9a3PcZESQyfmpa00S8HVDaPXbN
GoKqr7Yqy2iSHDVxggs4S6IDzppTIo5OR0VHLQHvSHNefvpcPpfTmJZxSu0COeeE
DvGkdoahuufv36DEXGpYipzS5kIpUQn9oXuGVXETq6MQz5kk8viPB21K4wN337BV
Ul3J4COMDCs79dXjyQk02KDQl4d7YoRqdI4qkYjiZNyu/QU6vnybAQGc1MOeiucd
BG+QMWUpr3l6enRo2cc2oyU6lcfOvyANOLgqxb3qx6X39aGMlnJdvKGtoPZ660eb
tqoy909UW2yLuxC39RXQaJ+4dAvwbTockDWtteACfACTQL/HDCoKwqxwfhJH7bB3
UDzCKr7UPyjad5yT/2yaciFofl9XqeuNUaSZwYUgLzy6qApfdrjy/WN9xFRCsAeE
4Iws0YkyuozEcGe9WwC+hCNwHAXd62l9ZnPkmSteWWjMwpXzHnJ59O4mQBThhraS
/cozw/OGdJaVQg6vxoDXnHm2uVCna4YBJzBmLdvWLdl/ksmbykn0byYbGYZN0sUm
6/UcJBTVndtgt3H3njGtA8rZsOKUSoJU3noV5N1CUf/nEXCPE6/BMkMMKjd1WDmE
o93pgfA+kBjx1zwNKZKra7FvJH51QFn6phhb0GPWp26eL6CAbIvgYIQSwU9wnAB1
WrnStXRYIAZpE/7VOv3OtegyZnEkwq9D2pSDdrSN9IFWEgQiuFVYhL1zp8PrNiJQ
xp3ods2EzxKoDqzOcoUR/fSAxMFy3GObJjUIh+2MaNjylCptE+V4flua13y72M38
xkI7U6KnQg3gZVMq3Z7k32e4miBKB/7dugZE11hMm6PGJp+9gi7w5jIWzyhBuBUS
8F7Ib8pKDDrDEMwnZOOcTDpf9qndayCSQ+Pi47VTSzKoVlf2qKFuEAMK99hum+lV
VV0QFiKBnMwz813ZQ5ZHkveaf6mJloaZFCROvvv+Bq8JHUjHa376A9z8dMDULb5B
2j6P3u3Fa/C5CbWiDawmEBj78T/XT+KWHE2kS7hUKmacIRKufVY8JbnleDMIxpgG
GjN1o7FeKrtJSMNi/4uxO4Wx9LAKMjOUlQu4zU+aCx6uR6ZCK7ZFPVdy6TXrpaCQ
w6vOR8ZxBSsNBmBG/z4EnAZ2VlgFO4QpuJgA9ydrkxlChVSBxaOuiF3R8WSq7vlp
ED0U7hPi2VsC4qg2bdw4YbmPUJeh0sthDbYUnToFcQfu/LTSQtl8PIlNp9dDn2cZ
6e0WHiIWOR6w1TSS7TW40LWdh17R+6Diki4UBBsRZ655WJBl1pUsRRcVkl4f1EE+
aygWnlnPp3pWy3ZEdmLW2WKQfDnpvzVie4xHLa5sLMWWxCEZlmSSYSycTCBsGXC/
+vkaVke59EhzNJCXLI2zXlTILgkpOAXsSCOq5So7dJibKiYMUkPVJ7QdMpFy56aZ
MRMV/wDdMyzqLkDsKpPoft+S03/RwdwLStvqgMqQRzyMRV/0f1Zl6cDbaHspDdgu
XMQZTqLABy3xBEcZAzWWbBiKbP7+xrHH2zfki3zJzSee6a7jayTArQ4diDhvMmLB
zkePGPNwLG+h5IBYrqq7CAEmUaHu2yo7KS2VIRt9h8L/z4I2ModZtX3GvnWLj2Iu
tNEMy2J7GUf6w/Sygnuj6RMs0eWsw9tMeZ0yhl2lS+yf6+fWJLiIaLe46hdQrS+u
EkTJsYaaKAZ+WjztFUikOHn7PiMdcPHGgNNkFrlci+8ptDhJuukJGinT5rqgEM0G
mZNAE9hFyG3bE4ISRmpFAA9j5xd99RKQYBfTgETOfE3bnqbTvPHQIdDww7JerSIi
A57q215+fMgAOif2pSbQZPAOuUZAYU97pz0O7eygEHnk8RIpskCl+M6aP4qH9oiq
FuZrmxZJ5NwtV1m1mTaqwQO1LVGnqiryaT2MnOq2J29UCgr1S5LpAWDByWOOavCU
SjEgxwQZJmmIeua7CgVuuka9b+K7Agkm7WwiQh40SdUtXotKOkQ/xBSGCVADogyX
8CvurKI6ygS6Ko6jK/QAqLM+3HjPtkO7Cs0VkNwxtl+cnK7ToJjfwuCQ+J0NaZw2
PDltSU9e/AGa7/ePbjlpDr/2fODwDYsZ7X5+fbyMbKcdB88Ye4CUvZaQ1M9TwcJN
AII/wJzj7qqd+s7fW9MevjZj5Jak7rzWosB+xc9v6sI0ZXWZg12KpXZt/nLHRrV2
kONfwGbMniZkeEMUmYKvBOAvSSe2Mlct3ij/WBfx+ThV8wdZGzlxY3cD7JJW8LPj
P4cedPgcgM0koenE/blKtfU0LVi1U6xLrqY6vlGLfuGUrZVa4E98sRcrnuDqFQzg
dhwQakmZDPZzY/QWfIHzxm42hSFsQRLZzDjQQHJj/zu7c5Bie6bWfuKa3yVUqUSx
VsB5NVvzy8+UjtLiDCJT28wQTEXkq2XmgolYq/qGMCrlfQKCN5qUBAIN4Cr4SMh3
A0IJ4IL+gxJqPl/+/89M/5jRUP0bG6LHIJpVUNoatB6VsVj216pZPERxa/0CgIkN
u8icMxpI/6fVvvXUIIcOgaKw4jWo8r39UFeB4X4kdD/mQDC4n0B/X0b7gq015fpG
3ZKQNa9tNSY2EV9bFRinZSSkUO7fccuhbJK56+ROHNnlrr4H3hDTKP9sjklaOJWG
79WENK+LKa8XTNLnFsBwR3u+ywuU392qED99B/bV0WrS17GhdJdTd0yhrJuia3Q/
Jaet8CWZhk87fyiebHc2dqLZop0UbNxi9lzezeT5Q2ICM0nsFfF4eoll+waupP9w
PfdIsbTMi4cTbbB/3iTL3nGIEE0KgYt2HcQnV8i7wAvgeCyC8TrAiWoksFDOpSNL
31Quu1kITGhzVwrn7DGDXbt+u+OMgFcbeoa5YT9tDTuXRalSceYczyjaIm0tRGra
yXHaF6GYHpJ4GM6ewPAVAo4cdPoL4UwK8xzvqFJINEmdN2jb8aN8pbJAvPI7Khej
fd+a25qMKxAWOW/IBxsX2F6xkvM8WEySNfMZyN+EuBR7/lXuVrrZEcbm+JG3N2H3
R+2Nztpn5LjEHpv1UHSu9y0DUPLKvcjzgpSCib7bcEB86fydigMh51wPw6qdqsHJ
6Zcf21ycP/veD2t35cgXU9c/m4Eo0vCn6wXzWzG70XBU1rB+qpCelkhVdGk+PzO5
uMqgJzU0vyf/7t9P4s+AErldSrmbba6rJ6uALdJtasG+Rw8rS09JOPU7oBXCzrmX
dbArrzUlETEHtFI6/EypVsP0fnyPUrWKVd81Idm4q2x8DCvjararJ32xfTUJC16w
vQ1cxkGo0wf89tyftuUJajvbdgX/YldIVql9nXST9m7OyoQRp05qyv4yjDBnzmj+
EwdNJs6uDkBQkHvPjh+2ulMTSQTtYSdOCM5/Px3YRXwDiM0I+a7L7XEqsTKZRLja
7xVRaVvJgjY6i/QPHajSxMvHXEq/Kn5YOlXIIpCyMKQ8mAjT/A3O477HO/8z7sIk
yaenar6C3MH9wR16HGnhr4pa7TWihJNENtUl/RiQWt3FLWelphZtaktEY7z/Kd8G
S0owNLBMtU/h5BBDRcJ9QREqRmOeSwqUVRVB2NGI1zfcTfiN4Lk9YrX9KKdF5CEM
KSjeM/clvR/IwmARdZfIjKdqxQlGGE0jhdmxMWL6SCpPiu88FUL52PLTHGwkzIGr
QnztEG6uXIrEKTL4d7jNoq9WoutNxKaquczfOOAHHG+5ipLFqRSNcIq03XI/TjTj
LZZVqvpayxRs8YCR20SNLKTMWD6opZEC/FTsczGmPONDEA4svWixZSjHMGWToowQ
pIa/94z1plOxCeVY/p5Q9XasvO4wii7VaJbTssgS5jNW7WuKt2bhMDvwWxnnWrt2
qXeTzdB6IFMjFcZyufWKP9HqTBPUY5TQaED6iupuswCw7PKLVAH0Nmgcv6tLanP4
/5NZOJ8x0APGDH7mO/hRcVTyS8s3EzyJEVzTDyOAz/GZBrAADEeaAg9I74wd3uLa
uUyBPoh5/A7I/xRCtyYbfns91o7OEFC3i7/KWokhYAQrB9r5qDugUjHFphmQ5lbr
LEcQQ+a8OFwktrs5bJ+2ltm0LE1w8cmefbtYTc5fsaEhCDwf78vR52AjOGOVVXJO
eCuPV9/fB+vL4rCEjjlWJtK4lLjdSq+EH8UAT8k2AcQtUuxbQeKvd62BwIPJrBPH
HNXTV8YMu0a13hT5AR55pmAJEYzoeOnqtjQTP+AlY4/W3wZs0kWM59lvehnEFg18
WmHsAxVVUuInbFq8xttV9HEfyy5HVYiHjAWwxN0HCBfQNBYZR9ekhumINtMAfInT
xo5B2aLbCln/NbHmEARt+Xj1xrZM3TNffQB+PAJ5KA+pT55kxtn/akgASKPfVs4h
mYTZW/7f5hzgzPkyhm4Vjg0yFnf5vUhxx2biwrQ5C0WjRD1/Q1o/PPm49mbja9W2
BfVnLsRPw/BTaRPflR3AnSfyrl4L8vHHpyZmv2EQuaAqmLgkkqobtHGFYYZ0g7Js
FNt4FuY6100I1yg/Sb1D+9QAHBMm8uFQPJ5j6Mhbg24fmGFPEciRzjdZlhE6dCpX
Nvr0Rm+sJ6uetydr5o6eA3ue8vb0OxkinI3IhNArWD5wEFVYc3PtTLECx9uoP+kU
joKKeiNHZhzSFsJhsF2NBqjhxQMIXrLdik9je6jIn6+gFK664LuiUaGSQKiKL+yr
5xkH9AjZiaYATd7LPXTa2bzas4RmXXU5Q5M1407SsE8jZ5kC0CvLDPZe/FzhuIhH
KrRABTYgwm+nQ+RqeZWYTz003qOcykgsizW2wWZdR09SAbUxBhBFQI4Uiz1Uw/Lu
SfuLnN0YiDVcXGnSVqyvuOnTB/qGTzlgR47C37TYKN9tcp8E/v8iz2yBpLxLtTJC
uDaEIFqzc5TllQ+Rx6GbKBMnc3rtx93y3AsQLVb5aFybyq37/wRUd3+L5ghIRJDs
9j0octO5dgOcrmO8s2OzlBnu/bWNnuxcExoE4mPq5fIaBKave6K7MA0R4gxLISCd
ssJEy8WAiWd4qQuUDe6WN+Kc3Mz/cNL+jajVoqbQup6QMwiqi0sbSGulfcKdU6Jp
cQFcGO5EqHxXCaPdl4TWcWsQiDSCLsqLrOjt3EqqioW/EoxAvwfW5NULawnudjrI
tfsSCFaxqcXckTKNfWgwdMTpVkPQWIhMfX4qvPDkQ5KjuoU7KRiKrrnOyGrx3r5Y
arSh7qpNSjPfgld+u9tau5rCu5PoW3RmXfdH7wrDfgrfUMwqdTcf3Y8Xjk6nnojb
XPX7Sn2bbocah1VEvuKwvJxuwi8jIiSluxw1HWb9yxNWTKGaVAA3xzPVT7mr4+Gv
85TIDqAW+Du9+2kf7E5C4wut2kaWgXKHfQIxE3Gr1MNrLMLG2ew2b3j2EMBYY5L5
eIhxYJ3K2uqrplQDG8dwNhNl8sVXv9/JxvUAf0y8JSi69wcNe0x8YkX6v+ind3OH
y+WMCVA1AFvve6x9NR2nVi1u2Nnsmb2+qIQ+4VZ91hb2bH18X0d1RUkorOdUkYF2
pw/1CbpQd/FXUxDq+EXWNFDzUwkMY988iqKmwIC15MZA8/uNUq0W4/K4L2gtiHPA
7wdZiinVL/Y7MJbLWJ61xFQNXVi3wAvQW/fXil6MFXVYd2ZY16x7UlGlKw0F5hSd
lbbJdSeMbMWNi4/aWckCF/DmjAha/uCezbXWCmX9nJD68gMmX8jor3xC1+qWYWZq
VRFTt+ocCeiHbw20Fh4dYs/2m7nsmqn1w0zlpmak9ZqbfyhtfHzhzCHsiiBSkGHy
bNrZMS3Qqgvub8JbFXU5kyDi0tnLP9iIxAEeURbrY0YEtKwzHFuvdsp2Z8fgLkMp
xfwBHvrhIZNE8CY21viPY8PBWQMsLdwiFN7edYmJLqPITMRK9uPPQbFHP7u8hpJI
ViWG2381XJedrBGPCI8rYiE8QlHgphFpP7pdjZwFVaZ9hxkFl8Iu7ZwKj1j6E0d8
28HFQWwS+RxRF3FqDp8cRsZnilquO5J4JfKPJ188NyvtVEzLMlxeuNpLi4oMpsG3
5ATwYZMq8+MFLfvYMSlAA9efJbcaF6H2YfzBM5wbZMYBwtkmbboz1gcwVPVRUgws
4L81VVR+S4Cii+nfgFKGg0zd8lYgNFrki4QDmDPMRiqEvDwJR5a0q51qGb6MZ9Cv
KTrrWb2BNw/Pbw7v2OdptmOI3wcuTFG9luIYlAOKv5h8N2ggN3l5LwxUecztQBuB
Jsqse1+7JZ7LKZyiJ+2HyIjGZrVmejh9p1/LJ3T1Nf3cFJ/UUbzPDxi/cGspyHwO
GnzK3kpXROrlDcL9c+82nGLxjFfn+l6Z8YD1Y9oOI9cMJLF7DFxjqv9083GH8l+o
XVK9SFWtPwquAaoMb4fXOwIGJNFVKSFEU3WzJvNkNmbM9xlUc34EPd6BtF9xcp5l
ncO6tZZahr//6NC7fMLv00dPLCrI2y3i4AX26deZxUBmgQX+NzaWmlRhEyMOhK/B
8p7R/bJYjOB8eXtj07j0ZeUk+KUKbTanvhUsS/E8/Gd0Rn90PrCJTDvkFjOnwluR
cpmO5t/tm3EJVfOtDIfBHA2Rjcsmsu6fZMsOXovkcpFUkH01kPxc7QmMsM0nLmVW
raFOgBIeA9VAmiwaMRUhXfAD5i6cF5Vtr9nnnsGHlvCg+FfQXII9VTWf4bDKhF2i
jf0uf8bWal7ihmXaoRG0LvaUMHdVbtzxU0hZYbYHycI36TggD1YMukSaeZZK5boA
3vi4ewVxrC3Gtra+RV1L7CvgkXwr2IvtXvHLriGpv2UOZs5PIbaA4etYUxGxtX6x
WnhHWsbk18RC6L6a6xWSOqHi4afbUi3sUNLxMtTWTHrg5OPClwyPUQxuHWJmF5BR
IILVIJkUvxrmJHwzSK+yp85Scvr5pGpD93U0YgE9K0pvHrTM7QmljYM76E0OKSgI
epBKDt+U4ILkJ65KjAPF0emBrR0+CaibW/yDhbF2J+d3QYxk520VwesnV8opVAy0
vtl63tFp/yWydqyNIe0joo2OvSjqPvvZSdGpJF65pvOM8mhttsb2yOnL8DJtltgi
eQ6i3nJCGHMsojc3NkZ5et21+aItvlVowRNFvrzn9Z/gbXVsS6l8+X4Aizz0A60L
bfFuhpXLV4n+SlttIeWMXnxZj+cZGw6dDxfHfVJEDtuPvvIhrJKd9fygEZoKd+re
N5iCDNhcOYEVXS1LvFgnUtG2BDkupSiOd+Miq0fWPgsQ9lWI6rAVj5cDCjwoa59m
XYTeWo4KH5f5pS6DvyUP3Bb1cY7sUzJLRgBzFJh6ZbJuNXhLVgA/Oqnjvoyqul6R
+yB8WI/5bEr1fqwR3rMSIzn7rqSkJNHn/nEdNpUBBQiwniroGQuY6AoP+xXZqxq0
PrhBqQvgabSpzxrnCr1ZDv8Ie6Dvxigi73Gd8sj36BgrCxJKdiTLGPJQ0pnKyzOA
k/g+k8kRaJvOzwoJQaLehk9m9QFgYy9HshUM5Hnu2UW4ZwpD5BXNIdMqXaPNAc7s
7QQ6T1LZ4k8Ys1XisT4BnFmOJQCt0r9S8Vo/MvRwXcRiyFrb/pcuooMkGya9QGI9
0s3WNjc9I8f+nbAPoVeSD1u77lKTlBwKK8gHey/4lhRNh8HMiVUH11NE4vf9AtIV
+uwsMMiFcMQ+dMLNt/c688XLQ2Lqxh8YLjZxxXBCzewlbbEWGDkMkW+ztmOs6jXS
AUx4FBDUcgARch4LjYcKeexccH2wzNIHuJoGsaYKNf1hjcz2lcnpcdpFixBSzFEQ
os8PKpVKcdO3qcd9sIfoCQ2ngMjGVs2yF70JzKATekQyoLY0UPPT4HND6JHUbAgb
bBSDZKeOBpkFXxglQUdKtSbVDFdhCJUdfSuetJo9sHaClMVM3iwUICvElMFvDVFY
7lE7+oshjPPrvgWFKI85wmpWUWAR4Px/UYLmdvSpIZ3u07i2G/tLLZHgYPXJoGNd
78RuMSQbeKNaSluhWLSWchBiKizOV19mcKNqc4m69cwcbKgxRvhNIVp5wu4Ryzwr
4dRCdPIqp15BB7aYtXSZzwWn4HTFhVsrfyjA3MZLq5NzNj1e2M6uB1sDhZ2N+hQp
LmxJfzPYZPn+Z+txXHZ8uTDu06k9UTFj2r8ngdsqCT6vowfUmce1xarJjPAtPuzr
WFS1LbCKqpmYLwfOQq8tWERYouZwGgnDMl8CLuj2Yv3S8Jd6KJAAhxmUUtaDPRQd
ewvLq3PgoYRtq6xyMUj+hXs40I8Oqa7BaO0At4i/gG/7/wQgq+v6eiHxWbWykypH
keE18ZANKR2JNv/ZRVB3pa6UGNWFTyUZD90UT48OjMHKVmsZKXkLRYuf8BBkhkhi
v3zjQUFDePHSQvxQid9cBNRbwFsiLHVrsH/j19WC++UlpOFWoVCbUWWxNutRt35n
qTkfTwmFGA+ls1PUokLjiEDpa7aICn+KsHEWRyCEGJI5+YkcRZKJj2zvzQYuGcsK
0Iogj1BjyLctEN02h6OM6OTB9pRGoZWM5SvA93KQdcOYJD2BCue672Dkkdbkk/4q
MoHyEO2MIVers0OWj1Z5kShwBu3uhJ9KVYNRFjX2+tk9He9UNPa0xjjlb3kwANEH
lB/NnqpiN+at1gcapbje/eNEuyrTgh/tBlYr0ED6QPaBP33VnScdZfRoOcTLfTZZ
vYUiWRH/YeVI/bJ4nhK5sb+b/37TjHgeRe7hoWejA1kjLwKJj+Z9jReUGE7NswT2
pEYNVSEi6w40iLBtgppdNELraxkKJV8wgLHmhkSWFQPsrmPOUIvgSugQw1+Xjihv
+t6xsZNoFd5Hs3O4lvLIv8BGBVAmcm/jrtHfhqW6ogmk5mAIOds1okSf1x+4EnSN
XL05y4GSafelE5QmK3zJo9vJrU99z2ZxJPe+UwdcYSIIi9C3WT3fljonTQoggjdw
5Qh7sJKJBAuvGXDMHaUBTHOH9+TyKR2RqvieCgmX8cwuPgd2Ng2kc4oQmKFCUfug
QHRVH6t9i7hG+J5uLwNCX1GAQufcnPB85aE3IT/Ttcpv3HRbKwc4qd1gPPo3LTxe
x/8OMnLtNmTo5twUmB7Gh0g8/KFnTwLUgsawrUk5ZKyVI1hizRtsVoBvFsTYANeQ
G/LOClELGa55Md1MO0/+eQUHLXlGAKDKJCVRVTXfB3aBPfOt0l2KOK5pmNiwmGBm
0arL5/Jk2h/0vl0TORA6rLONrbuYwngrQlN56l5mtEd66hogmRgH8Af58RSvW+qY
hHRzjMgGBLMhviomrjQlrSfB3lx/5qdnfHs/0cN8Jnk+9FHj6qGsrn2lbzqgr3bY
/u3ZZI6BcVLWO8iMwktRUKK+WGw3TZeVfW5wkzgqgwOtNETWdYypgh1hNRffuz28
KtgEWWtncxKqpy1f6P1ZrTxirF1xoL/f7QGQVqHUfr3n2aUC88iZCugSQLqZD5Tq
iHnlksuKfYoyfZ4tjpoWK1gAW1cL01lGiOfTsa/lHMes1UkRt7kAfVReNf34P8dm
RvyiB5YwL8uSoCIEymkTyhNWkhfzm5YkVru9WiJ/4zgmOZepaR1LYdbMzcl1iqtn
HX6x1UN5NmFfvI6eiw6hJwvcvHiR1x6IjR0gJC9d9yi8Qfu2xKJrmntTm7sOcWSV
WYgaxPRwSMwc/Ax174APtDrqrU8Vs188IWbXaR913+qwd4I/VoRDcEyW9fONRFNK
5MSE1NrGqyaD02zclN2ugp5K1KofkfHtYsgMtHPR2OMlDrV7Ove0CP2H+XN8c9c8
w6B6j8kOH8F6TucIOuxzXjBTjBi/9SD3bmnn1hpg2ggEBR9LAEtgAVW3pmFBgFAa
CXF3tl4hPpP4G/mOAm6nvgMA17kkOcfyXIiZvZ8H30bymQyR6zYFQgNemvafSPNo
1MZDm9Q+oU+7YuehW1pwTvRNmNkLo8/0Kv+eBlHVCWhy5YdxqAHAcnwvSzN7W4ed
4myOwqHDqNGmHo4NvK21/327pzpw9D+zwq/PxUMFbWcF3IVu7ddZQD2ne0oMpEna
i2lw+Eu5BGJ/6GoYCCCsOo2RXy+UqcdtaVgA0Gf2eEQrdgn/TMgebjkc2QEAi5dU
3aaY5VH3KElPNia2mBCe1tFaU/KEafjT6j4NoWnqZTxMxRqaSQlfhUYPWV6YgL/a
zUJUZGFAuql63C4VD0KkpoacH4Z9PuP8vdU/wfNyxdh3xN3z6+CmCFY4fgXtLzmS
s0hGV4M+TOE56ERFdmDQr/LXNhLDHgGByUlRJQIHh9Fw7JbYflkTjuyDtLThw7Nc
VXjPmMLQ3enDxRZ5ZwccNoXb8Z9L3lMkhE4z9TRJ/vPtfLBk+Qn2k2YJaFd2LooS
k9+vcIYEUs11dIlVUTH0ltlEC3pXYXwKpFdIiyHnnHVEt4FWM4fjmXEgGBh/zlSD
ssVKgXq3D8XIgCEmEf6qjSIezoTTAUBZrhM8dSHe8lPt0U0tmLM6zJgUJeCqCPWk
s8Lm+rDp4KpnZ4kLGmEh4qMeMOiFBRkmBSfCFMSQeJNKKSeVU4gcU0OM19LxjyTd
57MIwf4Vzy7mpCgofZj4vNvm2T5yuJdVaQQvzJ6zTVOzBQqAQuI/yRl2pJNO+OQg
A0+vVIBuO+Qcw6pIReNyquD//ESVHuiEdlGXjYtqHhjX2R9h3Qtl7ix2MVFKx5K2
lAQJ781EKCIpBJ7FE9Q4FPhZV0qBwXzbt3WiKbygHtoODbPz7UlpKY3EB4jbbCUG
FoQpKmd1AAzkPksD5bCLOpq12f6kDpdhHRR2j7aNUJb4fxFn+Pf0LzqhdFsrBNcK
Fc0Y/1xoGb21oUe622TMxmQiyMXTFU4bK+qgknY2SDYfM+o4zbn3oL8zboPsXL2x
gcZV1eosVYNUhDda19YZi26DFc/3DP3uwdRbcTHXihcdxPAx2a3OJVVUMo/yu2ay
geJcGb3hCn3SyBL0zYwya5LLAFygt6/QgljqXYLnJensC+tXwXTlmsPNnMDwZd/S
R32uL8KCCXcpuBQzlCoOgUP4iDxyy3s8ZjQSo2Xrt4ViL5HSrtPO+rjJPvQY9WIy
0EeZiemilD9UUM8zCe/mBfgjoPu0dsqMPCB75MSXexuo1B1cbiDvj4ZGACjw54p3
oKK2HydtHWOMY87qDTgG2t5itBZt8Le2yEXuJHBmsJ7ihHfvAuGmm5ia/TPzZBXn
A12VScWZ14NmVfcjyD4YRbOBlEoVASute8tC52+RfNpAD2eSMeUM7gtvHN/r7SbZ
r3eGRWZfKsmmpyFaSJjH00jAPLRpfyWm+gRa13EGQDQRvnhf5nZL8H6+ow36d/2s
yz7aMSMYBG/7NwH2BtZNlObbgRHWpfdDc8v0tUBl2MOcVNIOGE/MmtDim0Xr6KQE
bsDD+mgn6fEhmxP1y/RuB6pg2i8vSk4H5rusCjWkAvBNMPF6vXEFVST+cBnuNotO
i4zmNJcXscBdsWedsODmOvsd8d7du/7aa3rLZqZJpamYV2bYGCjsV+KGLfxRy+mc
G1w2Q+4nn0UopVlRjZObXJqYJ8RFITczRA6S2EX6E9HjTf9yDBVuFvTWQ9V3ao9y
P7r568ev+J1pJegpnyKolygEe7dz8Ir9te2K7lqqshG5CkyUEHEz2oqM9LdU1meV
c/8YBlSPGQ98WUIe9E6wqJTYTviDQUv2/ub9gmJmo3cl7+3QaxzWq/wttCfhXR3b
PVyYO5ATEzvErd+eXRtHym8GdL21OgP1AueHMfsD9eWGLzR10Llo64o1SbfBfL/4
8VmPWMbi01NHnTUcyOeAKehbbAMIqjquXF0ZVN1q8U0F6U5AvGC9JqP59A1qmENB
fZ8RcAw0uiSwiBj9/fKrWp0om9BaZNNa9pBvIOwHcP7Lgx5f4a1LYYsVff0K2vVd
q+d2pdW9wq0/poOXDZ76z7AwmeWexpbosRZK05F/rRfqY9Yj62wV22VRWxmVZkM/
8OOZsvPQeu2cdlwfU6H6ueqxK5itRf9vxT2jIJmwRcrLcZTCXuVfgrpUJoxWjIni
j5U3Lx2ro0sxNqZSfCPERkUfHvGhmT6PO0dMTFTy7OydnLnIKKD4ZMbAdHWBEk8C
eCRZJiX/YQtSy6CgXbMoPOUA5y1Y6CcAZV1M5ejK+hPCmdB/ALO+D8hxyPexmEg2
avFx9K+CmPRw8ONdY6QXpSN9hRtwuIfUAP1njfkqElv1ny8UFBh31thsDtcodpls
TgTd+LKIznM2tuTGdzcXB1pfsSKR3UjB80A6/y85xNtYcFUtJG2raup1yVAMebdl
MT4Ob/ZQ0IMVMYTJgRNMNmolHuU0b0yyh9JU1KOvW79YPjU8KJFbDepB17CHfrHw
+Iki753q2lyeGPO3jNG8f0RTPLrM7J6TK4hWMA8n3djWrnHUfMjW353DrdVBYZRg
nMOyAbb5oMvfKFNJsrTkTMpL95m/Ybu6cVGSLizZ5Z80yR2oBj1z53MeF6ABZRRh
lvAuym+q2STAeXlUUSHpW++GGaBVT53MDTH+tFmiKzkNtxtvz+XAcdsm53R/O7hB
itka454dAIBC5z6kK12r7VoLdWLmCVhiwxrYVdITwnaoj4OkJU7ctyb0HW7wJMq2
T8j5U4hLLWi05fYQEL6JndbfGYELtmiBWioNz0OeJl5Q9Gn9FabHaFYDmzNu688B
oPyHXuCv13KTJQQMg6g+sPW5siIjAdpvf2e36iSGSibh2px51sZoPrNIoQNjrxFd
YqseQnUIuqzTKbYQ2NrSLo8R0BOeXxR8jxv9GNr5qenpKSODyqmWJEtk9hNmvMT4
2h086CsTrf0EmRkT+FTQVyuqGYczevhZCE1wHGLV77QI/94Jcqy/A0igDLs4Uwau
12nrzMEW2DmP8Vs31/hAMwQbr2iYaD7v+eGmlOy4DZXL443ndj8HUTG4kurY52Mo
VOXoa3ebk38XnVKrM96L+XmO//VzheGIYjiD9nwME9xnO8MAEr+of+W1VfLqg7C4
kPZJubXx4eZyJVxeWqhUld8rBCUYPVWe/g0mToBN0i/mB0i/Bp0NFFmTOtRFV5Qf
OhrANuCsIMBnZdoOuzjh5ee7F0RysDmspNzyWpEGgpploKcZI6dw3mMStz/ONSG/
7Ch2gujfCeZQM7NL4ptCuwPehqT6zPpYSkHZUwoG3WtHQ6rLbOnUO0W5l/i6D3VO
OHlxocVVAL5NB/s119Zt34InOpi391hcM85XYiXTL3xqdxrOtteQS2Iu/WHoUsWx
r/xvL1fVwakL2pjcWBbX96oIzoEmjQh0fZy1ij9bD+iUiln9/OtKg37K5hmxNNo/
9pacahwTh/Xb1osF661IP9X/b5nsgZtlhZ3mHcFAkMQtUJaFXccj5tg+gOFIDHR+
rbH0pFgXreURUCkilsuA6XCkuF99RRu+UvbFSJ1msLYoyZVdUGKrd7qIqnv0nlQT
M4UdA3+/6PAyyM1n7IIbaRFkvR8TAVJNj8Buhe6bTLibfKi8Q1aa2ZPMw0sRALDC
wFgPnSc2qJ9D5+2E+/AwbWprSVA2uyiLj0hWYUyMcurkfFMwwoNdoTMHqrMrlPGp
Ek+cD0okXwLX9CnEN/Qm5DumrwfVFSs4ikpTtGV4kxav5iFItIwmQcyEIoBfsLzh
slR+6wLZArtrjB4OlpkFRgfs7BzKprGFelbV7ky1UfqISgWABk8ns44odVjo+7Mu
xZ1y05WHHnt/odVMMdLOU+SMFp3Qu/ug/NqQk7TNWYhF/aq8f9K6rp4BYf4ZqPhq
XKTvLXx3VIT1sD/LW47wJMNdTIm7o3mPw2GOAVkl/ww5dJktE09KAr+5Pymyctl2
0Zkh35eEQNGW8Q4xbWUVVprWGL1/7GtSHIDClMOGJdlsrtHp7/SCy7JKK/ctmeix
7O0cGR3Z1UTT48fbttwfWBe+S7IOi2PvJ+uu8YQ58ZcnwmekY+ReNqcEPbwC8ywu
ji+OmZMBsWDZEAy05K48qCrFGMyhkVXFs/8J8ldPGY5vfTuqAMkIgZj46lppliWX
dMLxiruAK3RtkIIZ0xlnPDFryjJOX0BlFxs/pN+tjavFed1/UKUl+xiqctKuoSzB
138J6MuaMRSgonShQC9Q52LuKMxffVMcm3CygIelEJDMI1RDofr5WI+v4R9+xD9Q
fErKUtcPWmsvPX9Vmmk7DKTi8a6SCnfN2Bx5FBIt8aEQgeNxMAlGgbmHWyOXGNZA
CcYXS5x0xlCtmAW5YA4B+9ppOQ3F8ufrmV+wh9khYx+TNf/9PCOq6CuGWNjjaES6
z+rUV8xqC4Di/3vcF3f2W2IbF1nsbeeMkZxmpl2SAeKqeX+lg9PFfX9PGNWzqVnF
/4JUBU/ft6UvPlJoZW1cAdrAqCGFP/BL//ikykRXJq9XiYpNqhLhNYZlwWNhnOY+
B8TCOPtu9DkxcPtn4iFA5YSI8/IqAnMtXvLXnui9twaXG1bLWXah3sbmJUUoaJLR
eYqInZMPZWxvJTkFORoKizCrItiiKiPF+1kMahrTgH2nyL/bxPvBxgr0EHUU1tmQ
8o3uW85nEl9TkOkGzuYo8qffZay6oFwOaBSem4k/RcUwVMvLgjfbpA5iAnq8p2m4
Xi9kVjBk8yXLIQLxfSpWcIGU4S41UJWm+Dt/0vuyFYAxO0VB+zDTAYsWPvbmQUux
tn+Nc2kTDyk4A8eOZH1GvT76Lp7MZzTjIjOHY1P3/Y6CN4C/WJ7W/DXM2Qjhh8zO
SLqkMztkGgxQUdVM+bhSDehYCtAXUwUcPFl+n015LFFID/n/53d5SNQe0gUDES5L
/b9WAVVh+6ZNLgUL8V23jkP3+pRFj4alhGEiC/0F2hjwHBQbFc2iZL0I9CKfXCfY
IQqWilXCtrzagstBQHh4wQumkIYEUuatC6BPiqmqNwTClCIrb9OoQtvWpHVX4qe4
zbqkUxrdXHUuZKKrUYUuxHcJDAPGOrNNbIK2J5VyVdTgSp1DyKBQ+a7UMcSo+889
Ixfl04Lix+jRrmCJNRoDnxtaNzYUkY2mgReYQgoVaKox2sxOXF5mu0Q5OMA/o8Si
GBZAjVVIpboXy8euaTPm91G11JFy7xHHNsJZ9KLxFIbnwKy6jvG/HH7VUj0czXKw
/9shjCeO/Eb+VwsGd+e9Ud8g6VBEVp204qB7Akn+10SbwIMFFx8GUZx48H3+FWQB
dJkt/8ILP+NQa1xtoMs1pMEkcR7+YL9xUc1gbGCb/cQtQ/MeMqCgOF1OcDrJGO7a
Q9Si4Hfs2faIPPJLjthj5fonxSxH9gcROcznIeMoDpNbJd8jtSEzksIfZ4yVszld
SBu6DkcwIeCf2lmr2J8sLz3a93NxN8RLtYNiURcZI9zcY4WeV4v78eGbXESACebq
qH2YoIH0pqeF6bFZ0LJ7/JEs2cuhn68WX3rrZHYk/FdkjiOFXk50WQ3y1wsqW5Hf
UelutLeJugDBlQbONoYcgLeeaQMBZ1KDuWFvDMtRkKAILOUvtzPSB45fCcdaOvSX
MUSb8GKQC77kE3DVL41G3VXkFyv4DehiDBShLWWZVz7x8XjpF+6DmenTzELg1226
/UpKmfu8nuOqqE3kTZ7sTttDTgv8aLhiH5wXlZSFuED9aZdvwza1XHHSJTgrFeMj
YXk1QIboH6QkQPHZ3n06sr7vM8qw9aKG5Rbl8uSgh/c4FrHxbifEX2m8Ys7+SJa+
0sTeb2ZtwEcSNZcpz37gSWC3cFA58MZ8IIAr1IZRumT/bWOEvCo2ZiJTjRUWVhk8
/HyK+L9Bqg0/CnZ5WaV/O3TV0BSbKGzpnGrqiE9NNSPZpaU3Ch4L6pm37cbh2tXh
eV/Ee4WuBjhfTF9vOQ2sd8FtOrDIfixo2LoawTwUkjswprF8H1hqqsCeiKR/YKDI
wbI5CHDLQi8R+QWpSsJXpip8LBL4tjYGTvFJV2vClDHp/MlUTp4AXxggimdVpOwA
XF8N2yUEHn/J7NmUuSDedHqIcVdf+0gjU61l63MD03OmY8ZdDQgkAvpyQAUZHUOp
19LFvaOPypGjvpfJoqhhk9pOocXNKxeaOQBqkuSUDSD9ySJcR1nLZBUZcuPDzZIX
Ja3hc4IUCOJiUM9Txw8g6Izl1rmvIdwv8p80W2OOJ2AFM4x/ggnfQSxFMjeq07Kj
FubR7zYVjHtaAFh1F5L0zpmAZZCo1lDL9xOyOAdzRGZh4g1fXKP6pDg47Yma22I8
klgW85TLbfytDRMriTVW7MrlVE3kSIfDtgmwHWOh5JsnV6cChSvWRdGKvHdmUu1s
X2y607gYMxJuVEunLMiCMq96arCv2l7EJGsNJUzn2dU7CxE4vwzykbXePAo9nIrX
/X2JxMh5WbYPXVPkoabUhVOotMPoPBrzdeetavx0ZP1WzQVG/bcxnYir9nl0GX3P
bMSRDG2ufa3Zo2BMo5zYNpheS0DBsacYGKe2wDFF3DYvX0esxDN7jY9UwIrqhm2s
tZLjwI3TK36w+tJ2dEvLq/BYFQFqI1Wzptlnbzo1vnPEl2St/6BNiSiulPME0VQW
mBOaXRMKfFn3aZG+kM5He4B5M1ETgTFM6LGhquBBJYAQ3TOg6Al8F/rtgC19SHDN
7PrzX7RhZkhryH73/ZY2A6uojurKwwKwwuAtWB1kGyeAiIBB9dkAxdg4F2w+bsHc
Dmt8bPn/5FRDfyhc4sFK6K2fWK7JRTnuWbLr8/jeu1q+SxzcXrGp7STUZlQydV9a
pL/ZSSjHBYoeFj+xdPZyXsTNEjn3ynvCkIVskm4CXV181OpaLSP4qobWTbRY7RM2
tI5Gq1b693mH5PrN6hWeQEDk3mqUzkxvRuOCaTwalEiXxMwBC4oK/+VkqUE8SMwC
x83WgGGK2Z5uqjblzPanMYJXSnc3eFwS2OMroTMXb7/9fFZOO+ObZRSY33KwT90r
gfCvkLxJ9qmIAAO9SkIh+Xvi7CTY+fzu69a0YUtcBVZNc/B4mLEaR7b/tiByClSA
MV7o3DxXZkzYf5NeGOx6EfoKzcQja3st9Oy88lqofvvfWBKaOE/fWkA3Ei4+v9j7
vY6852+5o0+GRPl4gtV2qoN/szuzVXl/kg8+GyGYfh0q1K2dSD049i9NQDnSnE7S
uPjXILhBmsRajFtpMdOCXOpjKnOKmsf73UmuwtKeW7Pce5YnOzABkoMvHLA5LnMr
Lf9ou3slWKzUG5E/rPrxVjFNOP2plzwoXowvfi0q8KjVFeKVDsDVu1deYucXpAVE
Wb+Qood+DvJxCbu+ZLaInf42qopaFgTDGH+w/+okh3l0dQv/LK6TQAK2DitfiGIX
WVDDpy3z6ixvrEniQ4uBEOv8B2dQ0Apa/VTj+rX/uKQ7KvtCNST9FiQzP/uJdb5S
ZsqueToMWKMVr+ykIyjjtd2TmOOHGaLUZA29zY5BHBrN2Qlw1CVgr5Q4Y2wbHTBI
BGObgPY4+6l0xBS43wnTcYjJ8064myKaqKNY4O6aieEhXgrTMhQ3tJ6wQUqFzxcy
Skzngbhnf6W4dYda8ERG4IOyRtvm9XJmI6Ry1gbJS+Mv46XQsty7Q6rnhvyByOT2
WdYPBWSp3u0n6r10i7R9HBRPUOWEbL6h7lPrO8/I37Gm7uQM3EILp2MT/dEkCPsV
2WH19Nx2hkcvszLnGKfjEyJ2e7GRNrE/QnMwgnpptdh2lnBun7PBmDZwHgA61W10
lVZZmopR4i8wsaqeq9wrsdX8p3gTOwwnQbOsXur2GIuIqjsHECk8wg+CGlC53xC1
MMF3qXNB8nQnGkQD8X+cRyvTg/uSHdoJMF9kNwE47p+b76nq69Ju7Nzugb3r+AzY
TXd8cbN0MVxhxQiFhwzdIrtMvVOZJsiF6pJkigIipLn/VLQHvW/Si4UUe4LgYw+s
2hZImrR6aTIVDyR8UAmdM632S+lWI6wCs+xFJ8/pBmoZVFyEPlcIJ52iy2ffHSdt
p2VvtT6OQeWl31YmTTCff/Mdf+oIALB3hIRTtTj4qGyatCh6Bfyo1xR5bas79Tik
JQnaZ5HKUAlz2J6nQRteRogpOQAP/n8OOGcSXESnxtZUxwa9l64nYY8nYwI9YCME
G66KrgrdkWPaVcMz/otXB2MQ3ezQz6tUuK/jyczPizaaZK78hSO6uyIB4Mtp0m8+
lVdltyYVwZ5+ntjU8atSWausP08uBX0N2kOJ/SdmWHQXei9DGfiQrqPY7/xZsAzV
o7zzz8gWSF+yi4b9yc5P25wzy7Kyvq6luL31C4T072fLO24pyRtHDRWPuCQrkoHd
m+XbTE3Rlw0wStPsvYkxJ3KucyyLzztIHsjSqIEV4/iLPiAy9GM1Dd3JsHvoynSZ
+10FjfMUb9rmLO25Kuj1REACWaeftDqlYUGRhyErvV9P5ONxNNi/tyhQm2pffr/D
p3Xr26kWgepDF/v6TIZNt3vzNwyhcZp3e2cwF2u5w9CD9IZFbFKf0eSFuHmnH+66
DsTKLCCJ+qQlFlQk9uRMs46YQ9Y/1T5BATKONZIn6xRRWrgPdVqVpQ0UeYCaBcmQ
IiSbueaF/LMf3Xb8IRnVKtNOlYyaIvSmLP5qG0VH55f9uOXXn5RVnjD1FyyatXIk
BWwCv6IX4fcOEXb28e4LGWJj6/ECK8m1X7sY6hxFYTKkgZSm8JpGjxyEd4fGJd9f
qB7jVw6xv6LXuxlQq/qMphQxPZYl+r9uGA7SuT6ggmqgyNM0hJhkCTeOxI4l+K1h
ziBRrstcQAXI7HDvyCB4/w9WEGAKJ0bbmasYAoLK7ZLzWNrXYHIWxgvoxBS/stYW
16Mku3B1gElwcXsjKUlx9lKF8F8iUoRwh2uXeKX6odfyEquBoIfzANyM0BeXWHd5
P9y/UmNDid05SXMzVyUsIRRdLYGMVC4aKkOo6viopL7+eDMiGS+sBnIGgRMaBTuK
ildzSdy4iOZJAvcFPrYbSqdKIq7BXOBOsVuXyMINRm0r935queM06fe4aIqaRrcs
3G8kOzpkMUUXPwXYjTDfAdyXj/MeaHgkHPZ8tLT6H5sB5ygMEt/S7Ge5BGrvlZnP
+f3qFi3nmK1Avekl0PUVYW5QoKrKrb4ksXvYkcwOpGHJ0mBFhEFe83vtejFTnAzZ
kiQgz+zFeDTKWrvUvBNvEc75ZQ0MKsf6Lfkf/oqcpqiImsQyKCZJm/F0IWv8OlqL
6m8z/Sis39VDMBFNKsUDWUbEvYWN7wNieGW6NKgVdFQv4Yaygj3HJyyfzCBQ4qhc
lOuspvFVgFsxEj1n17eu8dCd0luk7kdWKFNjGvDHMbQBqbU7eLJXuJHAyoXzxjEg
uY9QO2lZBktQf4OAdPA6amtJRlmbsT0Dr2PzHvwQv7kMI9fnJfSggUoIYvPPjzhw
NpT0q6zWBps5gHHY4SpmpvYwF0z04kRZ9MzvkW3KguMgqyQaWbyHE/6oo7VFTtLf
c21FjW7vXKd20uCebppZ1LjEL126/+FZAAVtfj+EPC36acLLaVWLb05Dw5CbqxxV
tzuNV/Yh6L3BMVfiJDlc+rJUw70HIjLCuzJvIvJhzv51jOqbkbw3kVTg3JB2llHk
J1tHyaBmmSw6vGpjIHeLAl6S371pAYMc1BXd7NVt1OMXGeCTkbHc2ffgXrcrK1G9
RzpVMtdnBeWatcWbS4c3J+MSCxl9OiSGzpX0a60ewsJr5CDK2jMg6cMcoHKD4fCN
3NU9EEzLKP0hu7O/nkdQv9c4TpoJ/7GtJwJbgJKZFNWSKS0O6ZfGsonM8pkGn+MH
RrttfkqFB3vfjj8CI6hdY+xcP9DxeR2uYXgpkedtTE2YKcqljGicq0L8tkSOaUlB
UcQ9XuYBK6Zcc5pfrWdiNIBtGErklbBr6OMLUBZRG3jaCL8wHx3rtTLYowEo9CXb
ZIl94ThUyntjvcZXinfmfSdYKI5dLLoqTjRHa5d0dLELYBIKXhUCX9AuUPNJy6pg
okkNAMfkZgjU+jr17LC+RWObImVPop15G9qvDfgLhWusaWY9iUdC7AsYUw0aKZVv
D/ivjTG9fMSy1b6/0r6eAwxHRjf2T4hSaLkqWNcv0SzZSiZgbGBnDhLWrQ/RwVxy
uROEhoIfXRcgs9Sr8enW7Iv7uIqmIsE/xIlDLixc581e/ND9m80k7F+ubJOfE6JV
u0S1XaOEXroc0suerMywXHaBauXHhWEjO6XNUClptgBKypP9sz8Nb1rqJLvvnz2T
zJbDGb76g5zQK9m9efHB72Z6i7+E9JU0vuCOdzTnXcXz9ny7Hagj+WAL5IumSpCx
C3CkIMSNRz1J0El/LI/eqxuJ3ipRqCGBrZTtcEImxPw+Zuz5oKNTxJmhNActFZXp
Yjy3x1LJA5DeKi0I/Nimi9ySQlePC7Ct2iE07omql4gxzwvmGKiLc80+ifE9OuVT
zzi4MDz6BJJiIaZkI9abah+eWUkpUBBJiPeZ8Afiy4+Z4KWDjrxNXqmhWy+4mEE4
9GUaU+jgyP7ll1nUU/9xjPgSPFLxyn0nZx9/GJoa+nUvOW0zdAP7saAVPF40Sdi1
Vle4x9WZnClqVbKp+T5FBInjj0cxNW1wxddwuAOz5kVVCRiU06IPokZ02r+iVH6M
rO3vwmyJDO8DqKPEtBDMOEaIBGTyM/pTa9zOQCl+vtJtXsjkr6XTBYqc0JWxCsvc
TZk4i0U6qcDLgLx8pnTCTSVE8MNuU8uqKm0z1AJGkFx4arP2HD0Y6TGh7YOEH720
YNNAYZ18Pl3+Kj61IAT9dd8WjBPDFTldrZ9IgFgF3lDHlHJ65r8z27NTpeuhOVA0
8PeCCeyF2yuD3k2ujem8/kCE4aPNf97GozJ2VmcMabvHGjkiX/A4fF8waFj4wQUT
TaJQ0y/Bh+Nf/9SLoOa/6M1pQs/IedkjBASuaOlNqeeMXEgIrYj1DGxdeVJq4iZE
QTl22t0RocZZlU3RSGqBbsEcbfWCQMPSlD8w3lpPg9i8le7TIjEuUwu+romI6TSI
zeO7SJGrWWIhCnTRvVChVUUDS+RlHepUR0XYpo4pJfw4yeQ1TA8rbEiBfJ3wie1+
uDXIqvI/c4VeeTGaLd/4G/QFe+BGZ8HJwkk5AQ8rJ6GWOtW3JvyEnTNNWTo7g74t
5duvCuYQDFeboa6rYRzAhQrRPvNLiTUnPHJ+mcKFMoYAsefXKD21uMXl6oCG11ct
1Wb3qlPfMYLqxZhNReOnqF73HAnQpZGrSWvfrGPW54pQcIWKMlxbDDM9TmdOCtsl
aMVI9qJXSi93mVplwtCl3czPWnEg3DWbEBeYnlqPcSuuYqFqfcC0iNNb63gAzoKb
dTqJesfnnJQNRqzs2yDiOaYQvW2wN7JBri1TUWczE9vJFDJr92EJahcWkI8mww22
1OGzs+BexvdkkbZGj9plE09oFf+w1GTcyR6wsJqcoF5fPWm5bGyICu+WrEGCGrgU
fWlVQ0kowr7LcKbSM3542C5gSrRegKS7keheTGo1cBVg+KJ2ta84lu1VnfnF4+DE
Mk0Td8IRbsemHET6CMjOUi3fttCilpzN6DqPn8/a0pyGdtC6jXi1zKrrS0hXZRDl
pJYdkFE7IXgPRsUJSKe3oAKfWoQcYJlkEm+STnhezZcQKdbYIx/onlkmx0qK7YbF
j5y/2YScV+kqvMgq/8Ft7TP9zKWF4PMGyXjm+nSo/7WafdNg6sllod/M8aWNrt/K
mtebir3l4EElkC4UcbRsPRvNU+G8/+vBfuR0vfaey8fqD5nOQRT/k/Vjgfbo5ngz
CqlFiSUSjaPKkTCjC6ZHfSD+vIRM9dtESPpe6x2mMklZOP7OFGXba3ZfCApQRCtc
cM/NfOIU0PQCIsYGOA2tFLsUHayQPqlB6KTmyfWpVP2WJs4J1FCCs6qozPB8dUE+
6F0XRFtl79zQKIgp8TnhKfRrWKybbmqZFEXsTH5sJtUqVB4Us29tAqtImbU+52iM
wmh3LqxecqeNYbwfM6T6HOdNcJ0rs5mutbxNybTPUic6wN5gIaylmy3cQZAxfpHz
d2GzTMWskE30zho0OSyZ/b/sNStfljFAAj7b4CGK1RHuv+kwWwljBNNc1VGG79Gn
UiSMx5Ljes/ZwIA6fBOWO64ZJEylle/p7eZ/Ks0WJ0v8jTrf3CKormro9/fvR/32
ItqFyKmlr/5JiHT0ScTu5gjhDLUX597A4HyvM9b8C8w1OUVSSaZsYvNrDYyM/D4C
Wuaf5rS4J8R22NvbvSEtKglP4P7a7avz53hGdz+RLJ5qrXLOymg8rBNltxIHNos5
Zavi0GJx0ESlJ6V7ZX8/YBotx2ZtdU1jeCqUx2csmneF5tvXJT7Ge/5dJdw/cp5v
As2791x+j25BQ4SL0+H7PrzjL1Rr9cRvFW6uAtdQkuLrz1XZzqV1i8AUJ0GvL8Fb
FRnkzGEZ27/LdR8FD3uYYOVVbaiFnAe7fC6RGXEx4Cju3QP2WPmMUGFmuFxPOiYy
4Z9AM9VqN/YShxDtH2R3TbdZ9EygJMZ6rdccg6HfQEqP3fuwUzPBC0zO0TaRYM+Z
awuAUFP3qnK8b/hX7KBWYv9QjMFHrwAp34C5bOYx+ySnq0fISSd4vqDqhGXtsCfM
dJZRe/Hdw+/JyoVG+j1gX1SK4/vGx/N5TexB+NjlndpXTN6XOvkNbU+jZuwV6Lcw
/ExEICwK+ISvpqhlS+iDmE2XGB8jVKkYGUSFhaHTBcoyiQEjAycc/1pzi+BCYd+K
eeHGf8k2yGY0bcq1nFC/amEhPV07sO0Zk9/6RoUNUw5Yb4HdFB3qTpJWSMwL6ha7
Iu1yAwXi/c7nJrKGUKseodMxDwDMhHqvDhflPRICH4je2/kC7bfBF/usoSByHw4h
L9jk+fnjIKF1YJkUNPr2neWeZNTFxBxaJnQiISXLoF7TTSug7u3sHGJ3rsDRLBnT
R5hfEz+VfK9o1IOvZU5JaywknkgtqX1IMIrVdf8Q03KYz3wdTDsu7cbx8hrmSUXJ
7w+GtAKBoS74lc7bjbebNi8G7jNn5k7yMiW2dTtx5FRQ+y24HqnJsRSqEZDlmRye
/StzNEOj3rXQI3Qg/B7sPob7RF0j0jaYizYL2xt7nHfUVC2VtDMB8Ajv2FScxAKb
MXLFJtMb5RMzPLK72D9Q3WhwBSnaULT52JoSMsFZKFzg1IrBGtehRdphC/dxGDXE
HnQ7o5Oh819tpAEwqDq7nm5aUbSZCoGCqcIaTUhxzQOICAqQSxJC/zgYiEdb9Whn
U9X0V3xbhDvMCsFxwHlAFOwdBN8gkFpPKUoZCithxWJuqvVjhkjIvc6w0X13YOHN
pSf0L37IILxCXgAZz1FCXxn/CpXEfd9my71WeJ+ms7bilFfEcIY4E2Y5AVdf4+HL
5reTv58tAsyQM73ygNQyrowhBlI5er98CLAMsqFuTfA3ncGXoI3jS8346yM/BuOF
IklJYG5f0gQgc+EgTDthn1/3+ZAZeTtV4aKRtdNTqVKA3R37GbZnmW6MbqY3Ge27
v6w1KgsB4mq9fn6AADKNKCsVXQgc2fTyasSYq92yCvJz2F1UZat/E83vKXkbHx9J
PDSrUMkgV190QwHwZPyEMQGso3+jSNhSFWGliJe1lfLkIVgbzS5V8ewSRREhNQYP
2ZmleE8Q+MsF8kEoRSKitMrCu6SI2RoFFaPfd+jNdu1O3NrK+0qZwgmEy8mGjjBe
3EUQAcqA8zrHKgs8+bdDu9AWMTcSl5SO1LSyyM++VtiaA4NPB/S7jhRJHsA733p2
vbNX8alfqolwczB6kB1+88ul5eR1bU+IANBsLE9D7buMx5bWjqEqc+yoQckQdEjW
maT32MjPXbBLYJhzu9mfeXmBHbL4Z1NuT8PT5jbE/PqDMLQSxY8mCC//WTnASQqv
qMDFRfepuqAZVpfkMibV7qPSMewDcJraBL3RhQ6s8EqJWD8P0f1HoQutoNQxD6ts
hz7GW5DzEtPDGMI3StwZkEaEPbW4H1WTWjYKPwA83QK00QvSwa1fyRXecduK9XGZ
inICEXt2jXY+D70X8x4LTPSE8AgtUsRTp+eP67m2MSmhf8ZUKDtLI7CKtndA3BIr
FWUASp294Onx/j/u4QYlc4SNi8BAUhnPGXUTgemqYRyzBOJO7XImchPb8SHtO+KA
KVpi2j2QkxZxOM/rYicX2/2WNCl8r3Ozozq+dL15IDAE/RSzDSmi4VTcFSN/1shL
VrgdErRm2dZQ/d/mMmXiDQLmnD2awEWOwSBxFzEe/TXrHrIqg6K/4eWhDo3vV5rd
dly2Ha49/tTiPDufyId0sH38EYtCVzndCE8hBMsMP7uDn+36mPpL9SJYOyAhtzRW
/UzOptKx/MwlLNPbk4w1/Bb4+KoYrXBvRxh5PlplmSANuFLh41QY8YIl2vgA00G9
xmGYBkdsTHM88s5dmm/KjFSIWX7Ww95t6/VRC7cjk2Oe4bnqN9BJVle+K5CFdV8b
Sr5Vj4VOk39G2eChtvbOjd8bQw5Cj4VKucVwJdTljPq1nEve2DKWxoYtkX1JzVDr
SadW9L77aWBP/6+u1HBPKx0pi0t7lmA7BYDtXfMNuj8wAKVLpUqgQdcuFkJY7bLu
uAeHtvoYXr/OtZDAYBwRndYLx+BLLsAlRb/dbwRoUuyqqLho78SQlOrzQP7w9m2B
gp7j9FqO8joBl7eMBh+bcfH07uaRJZx4fiHjWAXyqzo0szpP+T1INHjh+2KDfBLA
hA6Ux7ySIoEFE+2GtDbM9nXgV3wL5JMpEjIEgulI2K6N2p9Z6KmjWtkr7YZxSEcN
3/1YdvWIcSAHPwJizES6Cru+S9KcIbqyQBOXGSlkuxGqB2emgCoIVCoEVxQpTWOr
Oka6PPcyI0jQuzrwtNUcTFFp+T/D6HjTAExoiPmIGhHUWYlOZZPSfQfYCx28L+YC
oEFa3897tRJvJzyDTur/Tc+2RnjnYdUFA8oowUeDhZ3r50hhbMe/asxgHlKUsnAg
/XNKQml4RfF6u26QUwWhNocOrh4Oh1WCpVdWZScrSurU1kwLk7PlqUsGB4/XX66n
lShPh/vEdEYfJ6KMWIcCH7UDgIN50o47Dim7C1d+hNMX0Gls5OM1BITnj6k9lq5U
DmFFb+vWkNRohlRvvhlSZiEh7m7FmtpnyxFgBwEughIWMzsp/hYpkfPw/Grg4Ia0
AoNCN/tAEUyt5bHiy9Qhp3Ek2y0SbR00rtDjVbM2NkpYI1cE6nkZoH2bmzyG1VV7
E0oaTJGoSigw2M+QNXeNFuf8FggLUP/TIdiDAhpcDPEYkNKEhWm8CGUcJvhkgEBq
oeQu9oM6HpcOFN3K25pMAHWhG7Zf6segScWE5zNycTUFWYA3ceiKX6EN8O0uoKOp
yjPO88DD4bpS9DUclRIvEQWyklilr2jEvqT+O6IAGR5Ub3kyS9qfmla4J1aAsQDQ
pZFuenIk5a3HzcO8dqNYmUnuMWUNgSQ5yc+3wCWr1Wh7zP/qGbToWJa2yIW7JBMG
i+Mgd339uL9R1wVYlfiBnUOR1LBp+omiHSkNS9w5Vr2j9Ihf4yvS15h//C7qJv4+
6h0EbN8YwsimEqjMLEwWqFU5fMUhqd7de/bvCmMpZDiuxcM1EFrA+gFGGbGeUNP7
taiMfOW47tbolkjvDQtwd2reop+Njk+Glc9MxwTKBRGBR9pcZ2XFzUeK9q5TwkzN
QHV5JF+hsdxHHC02EEWCSCveyRVFhJFGKFV2i8kng5dLEsXQ5c2v6pe+MQwwd2Il
suuhxTATmswL29t6HhYRu4JdAYXtL/ZOjrW0BzDJUsVR6Gz4Q0TEfqIZ66UL/Qaj
/PjswMIETNpIuMI8rbggK9aAKUwQUnelSnDowjL+M80MaJgQceScyZFv76NCMvky
PW2O5p2H3GooZARM3Darv1DFEA8Njl9DhXHGtG+Vd9zi2g3nJf2N6MFEfLFdusFH
SEMc+p58PSIJSIwrtDSqBh4QAcbSQSwZmpvt0HIaXg2ZsGeS2fC97ZAMwXQLVFRf
lRwKXbApJViILUiPpjDJWLvcJUT5fh9oyWASXzaMIsODo2q/CHfwJ4x1pyo0QoKb
mHVC5QYW4wga/1lI7/ZbvGfTOmjH5BlYZKUupivEH9MO1bQzzm2c1PSslVHMFwfN
dAJnhwh7tnA4hhAODh90cJNnGBzOm9mzUePlreyXXdoiP2GL+9haTe6nIuv2dE+e
i3FcPeREoONq9vZJt1qjGPK5E8U7gfCW93BN2Bw+d5HwFhEEjVd0Tuo79+3UdKeO
Yz2/aJmcZczJ5Ugf2VuOct+2Ucb01MFvREqAKsGHMFVHmAV5dkQ2eV/rOPbbQie7
mWy2t8BXjXPBT5aEIHQm0/exUT9pp3ZagK7rOQNylgbbOZmUX2N2KKrDYvqaT/33
VivYxpYlcEjDDezf9dPY9mIDkUAqb1nAN7UkyHbriNXR4q/8MsXbSZvZOZY3IV/D
W4uFcdDeHaNeQMw+LsoX9/A1btc0nYfct8dsXdVxONPyL3igpefbfu3l2Irc2Zl8
ydLkjYXCsWOfbivj3+BI73nsYZuAaOVru0lf5YO5/jLUcsU7B4gKLS2ORz/Z0VhY
EhJ2J6K7baoNbHEceiZPbmX0sQpltQTLIJNSpQmdSAmd3ZJjcCwJO5ivh4SYSqJC
rG+SoQlvTr+aH+yKKUGKlsGOADiDr52iZa4lOuliIXroD949VbRQRn8y7qTnZLAk
HJj1jPm1U+gdrmHMasK68yYhXQqAJTbFez/nYPaCpa4vPZ+8OHjyzBKpprxpSvYx
LQA0gl45NhtboTXznPsYiEXQMwBXhPZynyrRcl+mGjnJCHpUlLu81tKOwKZV6+U3
EuZ5pO4pOjjMpktArr6Qd93mqQEQRb4wXxLYA7j4UAemEew30GS29iC12+o6xOOB
CEOPeIx473+bXdAaWRDUH3WPMv8AUFRqbtnRGcr27E23vkNIlA0FWnzh6qpId3Rh
3SzRukhk49NfZzDNSfqIu8eeeeFnaSvML6Sg2sGca1d1kRVnnU0OoZYtURNdcXvf
bzmAfTaQdLuX256DFG1rGJs5YIfVAg9v4GTfre8NkQ5wj/JtSls7X9MD0CLOzQvI
zTaRBWCqKUD0d4UaXKizPW9zsFUybQZ3A/3Uw64xc73Yof9Il1OJKgYcrt6hEIzw
UXIBrT/W7F5OCdiEqpeU52aOCjA/XQ0zE2ZpiPa+VRYYy6J4CN9JC2gGIF+8PdWX
NKvSx+5OsFgunIPrsUQXwuRN3ZSt+/FRSmsYBjK3d9Qw2eX54IQsAXQsDx7osCrU
9MTKkSgzq7+x6qVEWQOCyPGxjDfeNnj6iiQYqiOhW7jLWRfq1R9Qsuwc00y+hPPX
UJC0X9BbasUQ/Oa4o41ziBlNjli1wqUhklIRlS0E+JLhKOeJ7w0/lmuYv5Z1UXLD
dIH/81camuIyLb1jkuLGdYS0fyPIi6/Ag7fe/Ov49w505LTA7klKi8xoEg2a0YHT
FrBXcJJF0bnYoEH/OeTXZGY5JG7ArGg52RxXBck+s6LGwmvhZHNvX2XtFUdx7HOb
Hs4LsXo4e2Q6Jphak0xvc/ytMq5zYKIgn5PhZEEt3OBgGXdSGqwNP2CHGmkanHLG
tT9dmAdI6QFucKLvCzHZw7DhHu/aH+DuPnndWjCmeVWhMe5HgLcoXuRiPQvfH3yq
Kcat8S5u/4/10FR/PjNl3X+SBvHXGmnX3VV5XZFzLQPzct9ZIk7BnndOpJAU3P4V
pk+Yf50EYd+S0cHDQM04DDCoHXW4SdIgAvFiq65s87zpN7mzhy4aCTmC0jQHA0A/
x4qc+c37cwTIcXuQsiv2/eshfaKBfcYt8nx/TGd3Fp9ckd6vvKK1eBefHwuywyYd
dnBDTYgXKPQPl3zzGuFQldpY5NUpSqy2OtcxSsmX5EmmbHSnywFKDq1XwzhQWvjO
safZafs68ZloG9Rg6TEGxVwtzD/Y10qGOfu93cdtB95zyZpXkkDxvCPJcdDIegC1
oQYW3x0Kr8qtynOU1WlWJS06K2TDElE2UwpTTVXPizN/P03ix1X4uIsbLNi7y2Cr
E12EhY/290kScTqCBY7CIVu24V88YFZR2llqvVt2x+yNb7+UeiYDbGA1tW10ydyJ
hW6mkMdPN2FOvgwft4h4QLArEj8Fa7zM/S9GvHyF6uWDs36xeFnvLqiAuX1mduTr
sad6Wz9NKLqggYcrCG48nF9dtoNaarAYnSiWRDEOEy0o5WYJKLa0MwJ2yJsmhrJP
HzATJNC2EOrV/9vIKSfGAtiIuM6PQDb59iol5AF4afzxcvyhoVicK4TcPnYyCKf+
nHmokHbc4HeT8izL22TMGXTggitZ5c+j9d4zvM/l/O0GuoyIsna5cmQ4BovWtyeN
Q0NCIs3JfvKAuogW11cxvuO7cjou0+NdxshLJKj+433UX01OzprI023m0QrTJJZI
W3WvD7x18HzRlIGprBarjk7b/7ubC7E5UdvC11r8hfL6w7hJv+ciO35mj0qjs8XU
f8bs5zRHMkb2AkSUJgB5FGjoMdOVrzJ15UZWlWr6Af0fr8wZazmWe2GHQaAmtRKz
WH/RT4gin/asimL06cxTsFM+mpoqhoHhfXit4izGuGE1QCbF+fMQZhEyryZXUczb
Vjn6n8vBuAOPDqrZQU6BVMNgWwiOT/MbYY/YoQpIREnnMy4icTNqMCZtvu0OQFCr
IktDwuNiTC1HAefEd3OJ7oAHQhdtVSqjTomHPF5nfwdHyReWQe2ujHusgZGwxH+t
PJig9yU3XdKSGn9Yh4O4sGQrEjGoD2W1hwaTvDCKoBcaocs31boqK1ii2t2/l9Ls
00qDeLabCp06vNTW7UAX9T7atH5wUMBiicW8zatp/lRkREmcI/SzLTlb7fZO3TvQ
kTPqbIef6a9nDjJVh6vuufPpfHAAT/RR1IXjaEhVW+EFqFXDB8ackUNly+PvnkjJ
o2tS7H57uiwXG+VN936/W4sI24Lz9YmxQAVityY0dIps36K0Tpggfw/wqRkcHKNk
KjQ4vEyxxz8Uing2ot3GmQbc8h5iio/LDJ0irARaKahDj0FMsZDpAoco00xW6fqA
9RTNV1PbvbJVKrawarD++NBXD9Mx0gNMvowbGHBn3HsBAi2pImL5RtvW/VfQf+4y
fZHmBoYCUmIODQv8NQVUyAvhSgMJnXFCjiDtZ7k7H6tNRzPky+GpTLwPGQSGBJ+L
gJVhI/09PVZMJI7OVdjBSNX09Kb0RSDsfghCzRWmMOflai+iNGc/TDg9XfK7Lu6q
KnPdmI34IdHeBJZBCGgvje3D+GKpC7agAm9Uy3QJ2IsTnSmlqQKeTIj9CW3qWXtN
2u93M35o4l32j/Q5DHyrZNRC8Me29fQUNCLUJtSVWTLvL1kw5ex5qNtJyKWIblkO
vDGHMRi2GEHhCyas9E1X562UOC23skeSqatJSXaXPaNYxaPKE++6Ldx9xgGLSXxY
vV51ENOfp880sDw0aFWl0Lc3BGffqYWDNgx8IdPMeGoycj7lo4eo8vUJWadcZBOE
RT3OGSMb8QJmpW7CEUIDtKR8dljcheCP2hgmkqBbkYlrlYR3qJIlevdXP+IlDYqm
RYq3gCo8MvomFA4GEfNl/Xd3EnY1yBAseaPGIo/u2QDSTbMpq31Y8nmXXbXD6ka0
9Ph8pYYY9FueMNiZ35FKpokr/O95qPrkbMFNDn331ojLVI17AHnuk5dL+USw3xZ3
YoKWEUpYNoBPU3xbY+Br1pEw4i4U0tK+R2jyd3+DM+1XpiMFx9MeeawjP0ZsqzTu
ekLRjhJXtvYFpZxh+YiH6/ZLoK3EX7FkVCdQVpiH4ZQV1q1yVU/IugYAWRyWjQHn
YTGBGRd+9Icmbnn8er+45YMKl1N2WqJ7rAzFAUJDOLVarajLC0uRIbwm/CH5+nIy
B3ZQMye4pFXCFlEwYqSrbThiIDzLmDQYDrIq8v9/BucmSLZjmzr3NHMS/Tawd4wF
mF/f6BuJZ68kwNATUQqmTWAOVDpP3JlCepu7UULJdZWKMx9whB5W6P11xjZMFJnO
EVhNngGSOvMhQ3vPTelQCMJnEuxoEzTbvxGd4gmA90S5gNy6U/SYJVGPlDiGMt79
8MaUiovBI+DHtaSijtA/I60zV2n6Uy2mGnSVHXogvryvP7rLCWleOBAl2rhdqH1Z
SbPQWKGUPBuH1/Em3ZnlL7vrWHjbFoFuzBMN34L3Vw0ls3Ab4QXxPWyIjNtfnn5f
V73GmIx75Rdt7OU0a2OWhutxbk7PC8yutCTo1Uzbs5ECf3wOEQQHoIFmoYH1E8wg
qaNInnWj/6kDHUL2fza8pV0miehECCUs+t/VFXLZCdKsAZF1vGEfDkjLR2Fzayam
4FM4+EgJ7Xv6ppNLj18sOypMGVpDMtCsjyjTCCOjxpryb5fqzpWbm78YfosVHso1
aPmZkwmSh3tRmPFFpUkXcx1dmzvOAVjl/CUl6wiR+q3EhZPxy1j/j/V1VfzJrrVk
KfftwI59p3uEf7hW2NbS+KHS5NpNNQ4zkwm9/szzMaBMVcci7KnHjSzuOX+rpCcE
iIRm0jgzXlI5IyYLiH3i5WH6opgzw6uhIuHp2YcOsyPgQwDm40yrFVnSni/KQcK+
lc/en8cwu8AP3CelhrPTycnk6knp7zUwn4rrTamt4qeOuihfb7MFwwCXx1/W8vk7
EsJ/y8BHJtVA4/hKnVIymdNk4meZoY2c7gMXP6kCO7h5z4zuugyadgvzzgGHptL0
toLD/THSvQQ/YMONJ3w/T0/7lhmub2wzCV4pLC4Q8jiczjHkP74gK5PzygPxBMHC
NYFELsZI4HQoC26b4IEdYqyjpTMXGoMG6OhfVsZY3apMB4KMpLvAgghWCBiUqUEH
3GsTp2sftkbVtFrio9vdb0lqBmm7bWu63/eCx/01j88NBYPrCUguvXa2BtPNzPb3
Lz/y1FPJJMNthnQoHMCasacZTNZbEjbcBjs4OSr/ubvQhRHTssZUk1AV1BDYq54l
1XpnYspBCalUXKajYM13d29E/5tBEW98eu8sQ5oZLMdrAuH4DVOgOVCcDrGRgKIi
GH/nPj5cZdvf8CQ6rA6mFQGhwoGHL8Krl4M+8ONArylzR6IPl5fzSyloTZJNjito
DtzZsYMmyfFAMnoBi98XUvIKuh1+Hr83b2bokH1mSUbChOPkfxT6ebI/pzo8/Nqa
bvKkYXDCnjcuqWtQslBwQFUtPGU7UBP3YHGrY2gYyBb3226VhuoEohCSQCqItLFv
ZP0UrupyQZrsR9j3DfjLAKly7QTQjtFi9M1aCoXjjTl9ps6b3Bjxp1daLBfGUeS2
oSqY/9kSrtr4jJH/9BEg7RxfGDkxKqgsVTXCo6PsBriwHENAGN5UFZPJCLXr2TUz
iqlHhoElxqsBizXE1H6SFwcdybFOt9kTv4tBR+fwaKzy5bFg8oSo3Y1/Ng9E9O9s
pIybi7ezdr+712yW1NeHShgo75cr0hoeNJl7hY0QBFIWKPrwW1e1zth8+Up6y6xm
hv1pC/6iBzymjNYjEGwVBsRGOFEW//bQU4gpXuhMlr0HJrkjVSuJormFbT5OLnm2
eDREMb6ygczlWhVL90W5JpExaQ0DYGB0wGNomqDKRsRcHzY4fBLrujbkV3KuTlH2
BTZ1pOnC+chkaPX0n/3qhFRIMoaf2OveE/rmWvhQT7d+acbzrV8cvD2/HBuiU27g
N9+4C2HHwgPtbNPV9cpklnCYZdHK4oj9zaoosoXUugXj4tM10J66NH80DkL694fv
34xnihwmfgC+H52q55uKD3cKU+Kd2pDkHF7UPGTDxBJRmL10CUWMT8MgNMTiXQzI
Tz6HaVS/9aNJsV3ckkOY0BwKzWPT5oQLA8idIZi8m/hlMNCu7gXgPSgOkZriZ9+L
d9OkLKLGkYQSbMgj2sILs5e4RAMLZVHb0HX5c9qwdPaE7LZjZs55Vgir4qMZ69ZT
1RkpbZ3jazeLqgR1GXBh3CaHhQp3fPL4pm5QkiMK/csqOAtO2QkG+HLxVi7zlgyA
bHyS2qUmfDkinITZmPDOwyfuut004i12PFLg/lZYYhtfUWazu6peBnsWOrFBxqiM
G7F25r5QxfoyLdIF7baR1GQcvL1T8VxCUSVC7MdjB2popFMYSU6wP9zCWBDSelh9
C1Iet299ylQkCWsSLCx9HZ9QwBLLzeKYoI022s1fUoUyhYlnlfXk0xROgJ6DnzUh
FwrRPL01XwPxlddRCuBXUsx7D5XSOgSg96fEq2bhTR4em/68oYtfSNxD9FuIsZDL
jvn5IVwnkze1hiovY4Jqqvx1u5tkeIz54pZzqhHuqgOC5exYaJEv/+1pibth+LnU
edf91OK/XbZG1GOiMKfq8C8UplYviPPJn+u976iZjOvSVyCkaF181m2rqG7T7gMc
c1rcPkatDvVcj6UFwuFoJsVRryPmnX2oeBUDPlHxEkVNEiheUifQv6uNQQH52w6T
5/L72jrABDGkT6FZIdNTBPr74gJXR5inZj7s74CfUKoAwH9Yp9fC69IoGrK9/wcO
IpdteNf6F8o56Tmc9p4jVPoA+KgJ9c+on9TAHxjzutY/drJyCvdouHFI1q6j6wTp
YyWjOYzu7DBz/oJ1NEpfzJtyaigQJc6peTUsHqFnc9IcsF7+zTd7vUGIYOnfr5iE
yfjgEk3YiJUPPPNaiZcOVYawrwPEsX3aaH+Y/1OLj6XaexhlhvTQgDQek8SWyeyG
yiORGYpzKgp88/eq5tXBhehBYwAPXweIRWfLt2sX8DstrwVOlkw/pBiopyx7nsR2
wDAj9FX30Horgv1jxjwHW8pN1s98MoPar0UOpZgX99n3OGcLjzXdULJIA1HJGkUi
zlVsswIzcphL/qgl+9cDcrt4YPKC1fei6h1iYzQROmpMfgH4V+BVzPsmHLkdtXQU
mR7EhkWw1b6MiNDMgvJFurWaZl4UopOYwqRJR5Wlbvs8exyVoLtjDOEN9NKg7+1z
RuKOWq6V5BzbXDgbSFIhYjx4cr8YciV+bOH8y54zPwjb2KK0FfPySwvpBPfPXbm5
UVeuAoLhXgENy73E1kXfin7VJvhNFFbeWQB5Qhm7VmiDtzKVAD5v08wNBWg8dAJF
9Wu29a3e+8ozDE7S1ZqJsqo/kLF2vY/BlqboMlrCaCylIFfglkraWAR9jJaY9Mgd
ZBwr5Jji32DVkAINGDTDF2jYcJg9k3z1E0TDx0fzCAZBk+/Eh8OVXCwuTHt9lSfc
iPCV753Ugd7wgGodilrYIYtWJ6iKS5DQ9LzN1hqImWk3dkzy6wd1/nPs9RPF2axA
D89UNnWL2MVtpuVAXXU1tV1e29akR8OPM6/6RmgXXUy52CC9y41S+MlKpO32g4oR
N4X6e3yLc5l2qC/q9xTxzjeCwKITyLABNcmg1W4J4zrjx4YAmTrYF68ZUww+Ttk8
Sv1++JcvDofE4Q4yT5J6mjRS6vWvI4tB6F/1buyLIBhEH6KFW0EHfWEGRVXVW8yU
il5JQJaoUhqXoWUTtk89GJ62dIKBB9OCluOODMd9hO4ViptMJl6ko1b+HraAdEPp
BMeabUXl41jvd34fJG4l2y0MCfpJX5+g+q4oH4bvXXaiVuIm6Ho5eOFe2kiwfSX6
BNu5e4elnYvnGOxFu3UchhEKMhTr00ZAQkKYh0+sQz9MlS5b5lQt1EHnmKLiqHQE
zLqsIZZRWsHrmNcLwtihx9nDuX6ii5JJp/B4i2TuG3GYyhMqihDCPjQC54Fze9hy
OTe5Ula7rvyHf/WK/aCBeyPyDa2xAko/xp5TR307avCQyw0FpaAABb9MsCkP2F2G
8hgCj4UdM4MYIiBCZGxgxKf+lGwGvjlFh/EeNbtVZ0FNqbPaaeTdI6TxwVew3QSW
pIo7/xF8Jp8aYxpkzryYkjFRrad07KVN6O9g3slo/7HpKZaeyNWwXI+x1hZK/Tpy
BTWqlC4OHuHnvcw8VT4me7aP0IOCmPgSk+qhJzbGrT570VZlVF5L/i6BlWGzJ6+J
pZt7ieRvL+iTO1mlqWMpyRz6ccB+G+l6tKk2/uL4sSabGy8QOqY7kDXA9AhUZ+ZP
/6/mD9+H7TwjHi4b5GDsF1BIVsqzw9R7QmtbNVxhzBr2vlFcw5zdEa2wtIra5BEd
2yjx6wFKGqs86/+O06I5OGZ//6lCTF+pwKL5iwfy7dB595C7Obz1+2eFFWIpG7ih
V6Bx8Cp3qvEh+oWxyUd4g4N52gnwOmvbe4pPHFepbppYYOZYqFeeAEKdGPFlPpxV
9/Wplr8H7FzW3nBaq6OXBPFGY4Vbg3g0jxQZiGw/0GcJScrdHnHEcgQG77LWttFu
ax8C7sicjs7UkzNCHWzpwNMxKAYjJLrIGcLRms05BbUOGYvrCLBwpTL1qkW+6pwx
xYwLUSPo2ZLRkKYdENXSZIPY0Ogv7Kw9UFieNkLImKmvdjvYZJL99KkoGqgwXSrw
P2RPwcEf7amaH15x9yJSRLiJ6l30o9gz3Agvi2XYWpScmAvp+MIdIl/qWvlaFz0U
lYh0Ko3UFDhLEP1aS0kd6db1IUEIW6Vrw5ARlUImbAEFbDUl1AtwOaD+SueR9CAQ
OMJv0TQMZD6pxwjfF4KgwzXDkXNMBLJWx3XbgVwRb288eHDWumZThD6rmARllyL4
blmECMAbDRY5zvrzTU5Vdydv5HFcL7Wj3y5X7peC6BKMsL3tJWeITWTaU2cybosp
eTBTXwnVMv7y+g181q1BPHc74CatT6t23fYhHEyeOBsh+ATWOJM6Pm4sljPoo5W1
Mx+AEujmbDc4MwWnR7Tnm2ImwDbhKtqFEZWgrggzqwc9fIZmCiR8boBSsayqCMWF
RBhHYffjnfd3kU1/GfIXh2bL+CPJkatF5WAhdNMXSs/LVp9Swum6y5z8BQSebOd9
A9xRQ2RnhFhNque8BJr5Un+ohXiisfU+Ws5Zir67TBuR+I3BwFdRkdj6YR8IMbQN
zJAh3ya33Cmp/DOCQDWGJ7tkqFh2pnKrLsAUj/9Ro7DMnjoqRtKntn3i6hZsqZOq
lmMZ2JqLzrnjtxGNPkBx0+FZ0nLgPDezaJpnNCvCQkqZiAbXGqy5hQb/jaF4uJa1
h2aChO+l3ineQhxBlafc5qDlVHuv1W9x0GKud3KqKFjoNh97gDKxxkrv9nRj33uj
U8Q5YbdDu+Y2NZzH8Ff/hpWF9rW3+9c2lt90PLPxsCiwfT7pjGqT8HXXAhoz+GAf
MGuge36n0m1WK5gNw4BuD18e8nQaSrr1goKcy4oahc1u7X6GZSafz6NEA4pPARHG
fvrVeyUcHN6pgKn7h/tnMPo6XhA33L/DSMJIVU4cF/PsmSrzn219vAsIoVrGcuTz
YEq750f613I7jujOVDv47XjRZjxqDyY0aLLU2NYQacxnla6FoL9XS3wyEWGGYDBe
7FV/Y05Dev+IMyeRM0xto4lwRZjBS7w8aZKWmWAmj/o6iTHkxKsPNcbSMvZI/W6H
x2g9JNz2TPHu9uI8iAVWeAQepOywJ2svZl5iEAAgPoA/2Z8G83RKB7xbUVENa2jP
QFvYMTfo81JatrFyC5GvlPKX3LRi2QYabekPT7Pdco2mwvBfZQmWdXylHNvNa7gG
yeCsOG3drvw1Y+e4toGyjt/Htl+SfdYXr5uO1F73BgwD1ZWpIE2bhJvI5TmS2m2X
Kf0jUwKaLx3ZCaPKESeTk2dBVLl7tcTAR+Y4C/vU17YkFgx3PlGO7AHOcp4yeTh8
AkkMb/Ura11oE+JeVNpHO3+J6naXkHrYYiu4c5wStiJ+iKqVNOe0cB3oqAMtaKWd
efgAszyLv2lk+WQa5Pft04H45bwtmpkqam0H64c5E0BAHtyNjVIzqwa9glLXWYMq
G+QjsB67sdpaQwAA3sanNOHGpejWjopa+nT1Qg0pxIDu2kFJ9/7NXWQZEhYsykO5
C3p0pTfe2aOg9qpLSmR+EKvrHsru2yLwFBPnSSD1T6xuxpnNRLybIuDQp8SUF7CD
/5nQQWf/SUGU6GwOiWtLXvXVIC1dumDMYEmv0EPsrKBcx2FaHj7rewQNTN/oig6z
jsO5qn7PO1A38MJCNu+cCKeu7VwhShckHUcbr/gp/IwyR0BD0Qj5QmMxK1Faf9LD
i1aUMLbvbNydJuBAmNZ65yZE9jNbY/Z9mNo8Apo3PCX1UOeNb9jnkrHedQtVQgAe
bMdT93oN/HOVUo4G18aoZCJbE3HhKgGafxKtKf3FT4LvEiK1kTwh6mEcPnjJz+HR
B7g0G19rWAgjdp6/m4oQuxxnNrjf1EYwjYN2per9hAG8tYQ+el+rscuha10hpHVz
9sXwYu4RCioBxle97PPjusABVlAU94JKI9+ILgEa/DRuFzW9sVd025HoxPU/edkd
6SiraCcUd6yHyDyGLu9/Ut1SUikDHHqh9xyGIo8eUAGeCpjVC6rmoMzdPcfi7NRU
O0dkuwW7scBJ5T74nVpzZWVFhRAIv57s/evo3Lv3Pvzp6atuwa62QOug02x4+Jb4
mCLbwzYIPIO6MrX5riH1Nm6uTX4PXE410qA94Eo6bVv6QxRS1wYF5oq8Ux9k5JAy
owhyZrCxaDVTUIYsf62z4CQSngp4G5SG79NqO+ULHd74ZRIgACff8JeLTcTWVR4e
5pw3hRCGPnJSeqIV6gOmQhuQJWCgnP0jOp7GLUisGq67YjoeeP3y+xGJUUxcfzeA
cAB6TolMQ57WFeP75lw/oq2OfW4od2uuPbmcODkLw0qh5T2NKP08bO7bqtVOhpvF
DtNExjQNaodxT2x1IgVh4CG6TIqZ3jLaDEELKgthxAQHhn+QGwL/wFYTSJqo3YxJ
8Iqa4dR49h1Y+G6U8hs+UHXf47nglk4f2RYvQh4NMGENgmQ+mZynRS4WL/ItOt1y
YdaO6nKq9xSU2uPTSP69WxzIMmFHJ8lVbG/2nWAH4mwsdGZ5mjbJw0ZJqCJQto2x
CKWdYBzPzXuYh72JYewdc4GgF9qdpaBOzNmjfbNt41Np286xCumW8Ewe/BnasOaD
7zZKTlG0+erG/EKVPwYdwUKxl0thI+pUUKkb2g5q8X4WxAwAEwHCTKswJtY7BXB5
0Qc/8ZgGZRS+61yhp6xGf/vvAA8wgNGLcyeOQf9/KHdndqHVbHLjVwnL2Eu51MRp
xCfIqOpR6BA7j7rklCsPnZNwtxYrScAUBclRigdBi+zqpJU/jWm7mxfYHeRA22BV
GqJcPemzCNp43u3Ui582EK7Ylv9n5ehYzycKq0wSKNqGrTE6BsMIEPSlbopGnfad
mnJs9AhlU293n9VvIOWekaAynO8N/S63wjxwGJttiBVRYG2e0h2iRSIiW150Nswl
gb60+XuguaOHCGLXvpa+oXb+i2ZagFbElB09LBhXb/mqYQbL///tPdZnBI2rOsyI
D5KnBMbPlvOI1KKgDY0+wTkKtmqR1s4/Y7B8rhhB7G24FtpI8gHhmUkUwu2VjuKc
e5w/IHQcvXhIXezmIEauG5VGGlcNBZu+P92/X3Joz6FNb85TkvJwo6zFelvxkjBG
7BSeJ39H3B4aXrkVsAqIdM/MLJOgSRPlfH7byxkTCSf44V7OFwjXOagfy/f5OIq6
uIew7TluuWSZeOOvCCldQeG6+Kqroj/n1xxOGtZ1eaG9zYF0mReQjDLyBindFPI4
GL873ZhcLiPyLKWzzkb92vsUypl1LBUHMnTzCkqQyRlTCjc6FFuw9q4mbOuvLS5x
y4u/BZ4Mch5aiNbmT7OpzYpb/L0l9TKZ8OwuMjvokorLbFcefHqLfOqQPza/oQCD
IaSQBHr8VcHJGE1L9HWJcKIsvtryDkgwBMIavXrKxRsxzmzLhplgwqfgW+/PHCl7
0dO/jlDiV7G+n+MEg64tFsCenNqPnKwIPay0Th6xPDEJD6gdvsnEMM/nAsBHj6vx
0FvcuhDk+Nnd7ktVeKT84sJ33ZaS2vgbTxHn1Red8r9jtdIrqTAzn9SycpsXOBOm
M+gSPrCo6+cTHdSYHUY5xis1ZKZ/jNXaIlPypPPe+T83vn4rq1bv7ZBTeysfGebV
sbzMLq1/gG1i77dRvAtsyPTcSI9HgKRSWumHob6s86vXTmQrxd8fBwnWxFpkQaK0
OnR963o/EjZkm41v6TTk2HZkotZ5B0kwNWOEVao9bOI+h9dNrp0yZ6T2I7mqcSeZ
SYf4i2BRJQnK/LH0TKlybxvjBS261t0Je6JpDY5wodynfP2Cm9UiPIET6peB5qqv
yhjnr3FnEjrjHciLU2yR3nK4Wss48mF7iyR+TgI0qD8wEgDSGh1t6o590nrdiTRk
5dyvkAFa4u99fG5gYbRl45n00WzYxqxe/Gl/ii4hv6zSbx/9jGHC4W/CoEK6OdWo
sQKycX1FmeelDr1YtjfA0hSXxpTjL/gbqAKVp9sD8bcW0HBsYBRVnR6qH62WXq61
CksdDbbXcDRrffaP1wSwNYrkmR8WK0bmym2vkHywDBY7F0Y7Y5zpaEgtS+70TxBW
+vswFOTLh2eF9ZUz9Fm41Kkn8Oe5ZzYL6dvkD0FHmt3AdetZDanwWy4Urdt4sCis
DmefhzA2rFKz6BQyUjPJH9hyEvbcm2g43TEGv/NB8gFXzAqK6ARwwahBm4giGoIe
gCgocMpP4jGXDWFbqCYpkQHHqMOrG8NJTyFpsIuIFlOonJdq773QnLMm1gvddSCf
Lpts+E3ZV6I8DsYY4fOmlEmWW//CjHKnExFIEkkIwMOhlUaFqG/Xm+c0YsEaExWf
4EfZgYeIL+vY0HU+xKYujGfuwCTNY6X43lLppXg/26krZLcCsTY83xWi0qFzVpIx
5qC95qwrytwcCk7x1MeduD5tneSa6DIUOF7P3l1HucFg1T9QwtISHwyT/PcJIXkC
7TstP73rLYoyQyVQKuNYzavDzc2bjxeFlGDu2284TFHhe201WOpKHJ7DZ1t5CICR
RhvXWuV0WC0gG8gY1/2+3fcDbBWuhSw+AHxRQ7vNiXlZ5Hk4+lscvt1A29vpWZBn
H3Q9odlvS35zzO6J9e234Gk9ysD6KIlrd6rMglEoONAm7ZKKVAGezIIspNstY7jD
OtKBBHif9DrvoE+wlZmWvcJbZmovETWff9xGb3eQj03JeA/WHytUWOWDcTSUy5fx
KU/xtTDoi4hhZzokAdfFyMZ71pssleJCqOuVXgI7EpwP4SbLiG4NtiqFaBPN5S+T
+Dg/VhXOmlVT7VPioqDrXmORUHC1b6Oi+EmS5c0bxYBgzTMQeStVz5iZkuOCaCJr
t807GwmQvA0FPRCdfnMenQaXRyFccwBJ2Gr5xeVWuuC8GKuxKa7XSSZub0UAqhWe
4w5WFj46XZ6J6nuI7L9pbsW2Yd118ZH9/dSMjRZ1ibJWnc39ZgZ1VZdjomCMtrRM
nv8m0SgX1xlxpwNN+NMrl8zG73W3kIJzvl97Y/fFtM59rH7x3p2frXAXqj/UQdjn
236I0E3hMxUnxrwvOi/30WLX2aARlSZGRai2AKjXiP/ksywWuZVVePjvEyIprFsg
N7duE7PZ7XDDhHbkfI8w0NH/bUhuEL8ruOJQKMPfJRYZ0Tdv0lGdm3POjBRFLMMa
W9W0ME2L7Cw7/IZMDN8oOogrxjQ6UegyLhHK/0C/zvwm9bgvJvpbdkXxxEutw27C
Woox5LW6Ie2WfVYeIFUwI3UHLVMroMd7iDQ1dKP3YrdBAg6EaT+GZw1PqNH20TPA
iNMP6iueVIqnXb2vJA8TZ5IS7ztCND2N780bkPNOE9eqHjNmpRZsJ++81eYVTicy
B1W3QUJcYxbzt4u07xxjoS0SLvw6Cxvi2wMr25fl7mdMpnUWoJ6ZUyLgFsQpzrMo
V2IpIAxoWIrDt0y/rgGDu73MvZ6wBKkDtPDMi/uA80XswGFK5xsmC/HbFSizjNRH
u4gRKZqTTMKNfmc9jv1pR6aiWD9BK3ATb2YwQ+ChWWUz0M2LwNxSxJ/hjz9wP9mL
Z1eg+S4ghEbi5J+Sfinm6t9rbMwkYrbckq+nzgaODqa90InGy0XYjrK9CWBPLLYH
NE2NODACz0OAquKArps1r04liU0jDyDg7KUiHuJG13W7L8F0u3oKg28HiShwChpE
R4ukM25gxgzY62t0X3ncSJngMk7No+GTFKkLY2ebcZA8L8+PNNCHZNnASWyzr8VD
4UAAjklMqvV2b2TDuCnLGXoFutm8tvxOBfGEVV6ocWI8F0uCbvQYCqYlAHhvAUs4
Ckq6TR/2Q/MUN9JtHTldSZEUCbJG68D694lKr+xgRRoIgu+8T2ZVX8edNR3VXbN3
fgEQlTrVO+nfLTR2TWJZ+f9AIHzXlmJ5nPgBQyBKBhVVpKtWPUx4texZ8nw6ov96
u+QsUu8aMyaF6/v8zmQX20emUfUC753pLjdE9ESlj10BHKavXT768Zw2U9nMiC8s
WvUrgr8f0ZNsdaoJiqIxd66E92pCXIdoArKutZHAoIhUY35KOcC/gmI7UKCC15Rs
zDdONuGhPlyUe6D2nJhwQT+HgXjuf8uXjjrT08W3hzsLlHdJAXm/7DTn6W2wcDhH
UH2sx2DPGSlz/eZHWR/wMFN4wukEii4OlRs3XtqDHFgGqF1xdAl4Pkblvef6ZH45
/4+L5Z4fV25LBByB/lj67C5NyJjNXaj8G4rXKRpA9zZ6yZy6Y9mChagjxEE/zp8y
Mna7G4JLwSHB0uQtKwddYYs3oNP+nlmVCnhTurWxIIUWrJ1zKzVnszq9hYaPdAeD
Az/u5ryLakpzOeMNg4lGN/oRi5fLkCeeSTKDUobHXmz61TKERQGP3LCbAtcZ4e1f
vKflD80CeKuHs76ekHFda8tkjq+iuxb7q1324lHyvYRiwrV3PFjkg49BAG1eOK4+
dPDuFy8FIyGN/Qpy4SptPbQKzHZdx67sJj4zxYF7Spwr9G2ulXiMB1LD5afQOZa7
y+j5KYDyOwTKYQKpFihXLR9n2ZAUwhv981/zjWROjxUZMrurqwER5Bo8Cac/aOvc
jmlMKq/ZrIn9GRwecXYGMxf2BgRh56jMXnq4kktFTrJ9u2Dms8GNpEucCJYmxxjg
6EkUHMqA+49RlZ1oiqeR2YazU5/nKUWDdDMRS/D53y6QNVcuxeqltaxabh5zGto4
7XpDUnrDfZUuhRFKgallDUQAqOB6NxLEgzXsSPvALN9kTagGIalZwk026mqmjE39
GepknpVekuW5fILk6orewdCSKOTxLoysiihr+bWgojeuxtq6zTxoLhyarye0TsNL
9byIPQfwclezIcXfo93Otef6QMmmzin9TpNnvj+K2LBzQXlf2bFOd3thAUX3zrqz
syyBw//hT8bISVZ4T+yqIeZ/G8COtANSO2cPQd6so3DJaCGC3Q9hMB7tBsPOfEBE
ZWAUaJ+qmhzfJ9z4PgrYxCTcHMXftEb7NutmMlNOPolEjPAAmyP4fVZYY6fXui32
ysYSs5h3V5hX/rLhIywzjD6NOfw+bRPgH9R7wst74FP3iZfeQgLlsllEo0FwslKT
cazCRUTU8J3zd2Z8Ns8Qiq2FodAS1tpUeeWKsHmH530lVMPlYV2gTk8uBnyYm1gk
AME8a3B/kkYr72BQZs0+yUcv/OuUhaV9JhgNb5C0WLZc1i79hFoGeKDeKmhVvPqU
b2jQmyNbfGu4HA2PxFRaG4CZLAH8pwLmYwKVvboUGZW8rnTF77rqDHlXcEqVl0It
8Zi6VJ+KRiYB7nKojK24tJV8hEsxF62T4KTvcDBxs18UWBohBeOzgOz1ittz5LJo
tQwjFPggTIetPzSuYjll0X0dtF3wlHWr/JxSUiA84IooTJ7cssIMmN6jxAftLIDB
4Ior9uvQDtgO7PuKUm2Nva73vYk1fbyxk9BIrdSDBIj4HyZubX1meTwXYLIusJ90
GBBpQ3j3z001tMnpZM7qxZreV5U8WYt/T1VuJhRieBeQkHugJuGdyj2eOfQhcXEC
m5ZarE+aTJ0nQkn5YVZOxfyQRmtak6Pz+eVCCIGoCle+UyUj8rcSGL2jVUoXZr8i
8pamE7MlhpIyo97GecXqQqPIKVmGsGjIUTrpoUW0GT1y5YUGHH3ORSeV03Zbpo/i
U1QjkGo9+8s28kGhte46iJ7YKzKWJ+OxAgD1jG68BBNUC8vv5RiJqxq2qdBtoO2U
iRXQdfJml2V0ut/I/VDvCMKW+VYhBILISUuznjON6Fka5A2DYSwdRMkqRWsCSi68
RNl1O19rvBVp/RXQ+9a59CdcfCVesA/zPqrc+rhv9l58boL/GYcE72khjQsXQDoN
iwDGtUEKUWyxLZ89QR32QliSlSM8tNLwLXx7WZNJw5b8FvdMSPt3tvzfcwfgBJA8
9N3Oq4bVJN+7hV7tcpA1VHCVpklpCQHAY9D4hpvsUH4d2fswObejCJh39P11940w
Nprm8rDBU+m7URWZF3VbdiX5A9WHVxAdGoIlu3iquyZ8ppszDtc77l6h5UTq5+9B
xfZQaWt5sER2DBMZRMCpHAFS1vRaoD+2WmGkcqAYfvhY1G99ReFM2HP7OqdsgrMs
GDZHYPetzPwqOEls7bKSY5ZcvnlJODj0nCu64Dnab4bFGeCEvXaOuJvHUrWsMSBi
tc7MtryxoZ9FMIle05IaUO5l0QmJwGgvy8bpLuEog5V/gMStj3bO1QpzQBbo/qDu
T85RAERPDmHcktNPkaSkxL7fqmk0yLh7utXp/qqgf/PutBxiBz+L7bUNpH75VM9J
MYau6FiFM6Jnia1kux5rjg3RlpK1sCm+SjNJTpsBtv1MNwiAvn9s0I7FE2RXLp+I
7FDiGNDG3I3gkxxLkWEE7MhtP9oa1GZUBqqOfgc5eIjkX7U2a60YTnqjHRmFZHrm
v/8VStHuHYvjg7Iz5D+KujJcy3HZgwa18AFcWnkMoR8M4UohPBF3Eib9ta2VsKtR
1d41CLnP3xy0/dBc23NRxpxWPALtp7PlwT/7tIw/T1tZXt4aXBggGz4+QsTuPcM+
dRt14iHzqK22P0p2JQF9Q8xa80whiH3voib39Sa/mXjWlu6bFqkbF/KIgJwomavU
Y12VXO9Xu/ixM+P90IFdKgT2onXp5NehaMpw4jlyUtaAwZ5a0eO+VdTUcK1jH8TO
GwVfLsSggwRvdn+QT7WSDFViOn/iWg/cv02+SjpOm6uC8tJ5FptniYoQQeRvEJr+
1zx8/NXuUj5X/QWOKXhX1GFBEovsYEUX4V+XiDbycOvzXvSp8UMJ3ItN9KjolUHK
x572g7GlXCkZQZglggs5yfOKrm4NDn+/LpJ3p93cvtHmbdeEAkZOX6PvccS8WK4y
L5wBkWIsJqrQ7YjtxtFrSLF563sRklfpQkYqiJ/X71lT0dCRnXVr59+3kVDVvx7a
EsuQ7bXJEWlyK7e4QV5yaZKGJZpaJiFPbm61CeXFf8PPGRmO3lruUSpNAx7L3Zvv
c9iQ1m3ppUONpJS9L9vmKHP0SE3vk6jMlehWUSVnDIpTrPbjXC0zPPuGO5LMM0BQ
Vx/QLpsOqb9J720Oo8rJYgov0zp2plux30fWq0POcn2SgX2oZrsREmf6CW/WQdxU
oSzQvFGT+WnFvqvqPozOq/C1yv+jxI+XmMyxkTpGcHQJCFIEv62/yGjvUnS3FTHK
Zvnt5r0cQXf1PJrPiB7mfCxqtBB69lmPHBr1rRfZ+hTHL2CzklCg8Z2YQA8vDFg4
trKQrkDmdZA5OuHss8lI6PjdGVvAG62NvxhcqRIEa3V3+K2pWIq24ipTju3WkC5S
dWIThz3sFOd19N7oZQ8kuYOSRFrITALSn70a4arGDyPOau8d2ExAEeMVX0kfPMn9
dg2wjEpN9debay3oaEhSkG9/obRQx9yV4DNdYgIyzkdMvs5e+LqZ+oAWIJdhXOgS
pNXrl2RRoolgIjP5or2rU1i1vqp1KfjCgMGIe1j0Aol9X9+/YtranpJbnNVZkGXQ
jQlWd7hY4iKgSVkTj41ldB44X0qHrV8SmcLmrYtSXyu14o8TbThCRE+H6TuZDwme
BQ2O09b5EODCO1YehP7TA0klY3q9q562UHZaNFG/5WN1q5182jMCyHxYqyEcA95f
oSGV1ke7b7D2oSq7sdrmBIFEOxafPq2yzWE9gyiBo+YAUhqOE0Gonui/tAoy279j
KZkkipwAE11JRCVjy6zskGn6aFVE3TZgADfMiaobU2koy96ISaShJ1KNegWRa0aO
0SDPt3iq+8GlJG3UJY8dydR5xjBz3iKQT6BPlOAPb35yarH9tUrAK87LN1+DB1dZ
MsdQ2W78lkjjcV7mH6QXlovMe5Zfs/0NrGBxgyKu+acAjl+XPTM6akAINPg46AfF
2ioiqb0ZqzCIJVLUpXwtzSF+G3aOY/3/vVQNIgbYlmx6XkLyNBd05TWW71jxpN0T
lBKIKskCIS0z6idmG7g0Z/yEaiEXq5ezkrCBHQpcZB5EGi2iyCsolj+HdQkpq+lz
w7hXRZp5AcFSjOR1WVV5FYj9IeNBTqTonukgeRqe9Ufqf3B1i6/zQte9msyj3fdw
FQqu+4skTVAeWj9tBKWmI3xc7MH1ZRYgxg7BiV88/U04pNCjS8EomTfssNW5v8GY
dv6huxXLbPc23wkLBEgyEvivgV18SwWbnTNKMDHOr2900g6Mu8oq95QFoIf+z0yg
dTloZaHEiT7OyOChObWP4G4DtFaw3jq1bX8Kb0bBthRTVyMQ//184yd579C3UepM
RXXiTIUh2ER9N1vm/6QSwvOMoKa83pkS80gTqIZuICdPSbcIlvXJ9/bR8QgBgdyR
0oD7fyI4edrVrHbC1Nrl5W1onT00jDJy+cerZZeL78wCyMA96lTKxPfFxC9ey8dO
R/kWNvkSG0JdoehnTlDcyxvL1/hhI7xS1PHkP1tA4xahKVHOm2Aanjs0uENU/SPb
+nGopTgQ+qLibr5+EGH+iWcTNDPSrEzf71v4FQ+uw1PwUwn0hyPaELirq/niGAhS
UnvVv5Ady/aE1q/mrhCJtxn1ZTupzx7yjSxx0Ngpi4xWXJfwgnmj7D7+MXF06mjM
F/WyovS/DpUWyTurVCpv+mmsiqNfPwDqrn67B9LJCBiySJbLhUfoV4QUm/oBBgqt
78xcCm5fEpQ+q73qkTj6+oe0pgRvo5tV9t8nOixIAyyIUriViQB0hRrhhygHDR4Y
hvQ+qlSDu7zcd9J6pSs2OARY0J85V0UIzk2V+AZMa/ImLe2fMJqJyb8tIBhZH9EB
eSNT67kFlVZPoDYN5TDFyGn33SXN76tp4oiexM905RfF5Lrjn5sez38JZoO2KQLl
eLrNl/ey6j1j4zrSAR/bTTt+q6bSU/cr0I/MaNQF6TzGYs/5K4t4AeD+nG+9xQ6y
aKnklacoQt+RVqUZLRV2g/Cug2YlO+4Xlet4IbLxmEw0QcPZ8Ud5R6Rwu5sQS1V8
IMQfIrZx9gNiv9IaxMIkFFf35WmrGFVekgQoj4/ONjAWequQmiuH46RACytvtR/t
xbZkjzvI6g5PwNSKy10nMXkFr6l+ads2Eg00zBYC4+n9sSJud1hOvSjaIAm24G7I
LZuIwB//2dU3PgrJZ9OxerQizdTDkc8KoSToqPA0MNKKtJhuU5M7sfxAmGW91eY4
ReaVs2mGT7Iwpn7r2lMthJrxRoZXpVoAc7jqy4Vtuyo4ZnRDaf6VAQDyzqV93PV/
wqO4bob1dAiXHHMRi5pYrzPdZTxYCb40KoFrTnThb25Uz4Ue1/tJHmMkMHc9qkr2
rPsrGcQRqepS86cCXaRQ6lGiRKIGKLFsKdfYrCiD2E9hxhdP/REKZQItXIT3KCo2
Vp8KvYQ0b7R9S29nAKeK0WwC5WlQaMaEf4D/3xMXIxmpxov9pPxnwoiamN1pUcJr
CDC3PAKfbn32jmS3hsinTXaLZmF5pE93BPOwJmuwND/fQtQXD084n7OtAsLjATPe
EcayUg3GklltTZhKzoULdQRlAKiqJdYZ1V+F9KtJ0SBseYl8e7LmkCgA4fZ3Y/UM
8EFhpI4iPw5BR9wBG0csGIyqnx1bFpp0HmF8QGkM6N38jUAsrwdMwDj9COPYSLJ6
l/MqPrhL47SEaXHdQRXzwvV4TzyjeAv7h9svIkGfXfe8kAkHMpLOML1yADZ1YSmZ
Co20WaqD0lHgB6eYM0h3q74WTZEkfavRyr9vIZ80ku9lw3dGzYDYkWT2hudlGYJy
p74oJHh9YXSsW49uPyFIYSRyEbs+83eQDZJcCwFOlHfcmqA0PkALq2r0MaG+xt2D
7j79p3RyAH5r+DaHp2C/eqCI7E5mPibNlICnJGPJC/XBFkUnbWhRUevnWAovRw8Z
BV3PG8usz968KORtgTw0H2K8gA1R6qYSCyYs7JPK6P6EW4eSC9mrlgZ+FqprKdlh
Q3t73znYdUtuokj74H/+7VbRwj7fHZ8sqTw3ByviQcrW4dqmdsgbcMif3FPUjUVI
i2A0tEBky9ossA4aX/l07obrLvPezlr4lV8CXqTkkbQhEYszjXGO0nOIjbwZDkfY
yka5BfhEmRBvmOQ/eMVzV+SEoyN0x7yzvDXvef91vTSi8ngHXJytZfvMBxvkK4P9
/dW15yCTo5kFCXNmiBVA4wnGxsdYULxWQlJ170caRE2wzI0i02wG3mdp8bVFy/iH
/gJDdcaqegM/FGfuJTqVHo0vepDwMqmeLYZqVBjj+F3THaCN8jqSocXbHbCaLDee
HcwtCgDEY9NW7jPQxKGjuBn747s8A1gDGw9khzAS6xxIoNWkZV+KQSVo3mj/JVTT
HWvdimYlRtPGmA8D+/9u6Dwnl/NrIJP3WUToqz6Xgkwr78A4T7qEAMlCNdYSSklz
xFEX5Fa9DS/B+NFeEFxX9BvDe9/HVBnaQVWiF/Bsd6w4Tx0XQhULnl0bmK4zZ2oa
u0LgZ8wgN7bFiildG1W5f7Yk3IBHmvSfO/a5ByhwpyFMdABEyJJQ3ovVzKISY5YV
tMkx5a5n+uPRn6vrj5oCgzEUE7k+6UXhUgkqHiYI/NtQNZw6ALWft+R+Sc25/rQf
mQMKOmPVInoYFqNgKy8o0+zuDLgg4CpiOoLLB+jXtk2//D6qLnNq0ly4Ro1k9ee0
l02gb57FWZq4kQB0GH8tMACPDYMqtRqWWPzAkmXsRHTemCSCpUThQLfocf5S+te+
nuatQ5eCVFzetvRh9FJtgYnX/WxWVtH0h6D3w6zLHbHTrhgtdBxeqdNeF5DTrmiJ
w/vtyrh52NoVl7siMz+qReVL2B9qsJ+m6B11bTOed5XOFOosgCNh/7UwudLFVX2I
JDoSkxtHHuq6SVbvT3sMrRVJ5cb0yGReT0zd+RcCVUntOorvmT3eU8eKTCPCqJ5J
Wtz+w09IUB3vGEhLveSuk0iWv+3xzMUW/3zWU5lrIL8b/Zrp0Odt7sXnZ4pjrAhp
Kun9zw6aHBlg/voioNsRn3EzLquSQXn1QEoqEsNQQ6vdcP9Vvkq1BxMeeelPK1F3
7gtD4vSRRwdaOmkqxFIFB8xXzhDyZsfuGtyT+r4MeOHJSWmP4U0R3OG0K5qLmGvx
eyJRNyIRR1Vsy+2Q+hFFx/vNvsLz5Wyh1H5P4OYOTfx3HjftuUZdyxRhzLWv1knB
415KdCq33+ViLUYiPgCjnT1wCjcpsnJQlze0WNvr9SO6zqQRiyqm2MnVpZKLPL6d
roDcZWU6PDfZkNCl0Dl0AVUDlbuy5TwvF1ieQVufOPKHjFjUyOdjK8kq23z6jWAd
2Q6KymCmYq2dLhMJe8pepT31hndMlxwznsTWXc0sQKg3dmS+54Ky9OD7Bp8DjEGx
+Dnup/6BpWs0qcXBFsdmXhU610BxPo+Afc6x7guEhtDlwMe3+njnpROee3RWhrqE
cz62tegNdS54uWGsr5S3TiIn/0mvP75H0WleeVcL3iWFn5CpOBNKFUHMLqRoF8in
sLqrrojBUbY/Oeip4c5Ji8jjrwA55GknWeWL5LoAt0e3fXTYpWofU7eRo6gjEdX6
uhjF1tJeTrdoQUxDQs4g4Y5lI39DsO9FpgW1Rb5ZmBtKEs+zBXfkloc/XInkkwVR
hVi/KroxVlRwmtb4KS+yKPtcJr4Hvqg6vYdLjbkEdA+as45Ee2vK1+fgIbR+p8NJ
ilABJmO80fpUPJHF5QXf7mNopj9J4dZZpDa1D8tlebJ5krSWyx4/b59FFIwjucj7
kiSay3wj3eFXxyM494bYrIlo3+6M9wdf4TImJzmSzH6UeosKObY11uYuE7fdPm2w
ofqWjQiSlkRJiyoyit5h2BAcjSFpwltTc0FPFFMRKoGh0iFOKIhXu1WdLlUL9PF4
qE2I74GwrKTFe6X1QlClKywlA8L4RSpwEe5Qiczm5mANIMN0ztkDQSh3dDtqe47d
KsCkGvOuX5HB8X0hQAOLynLrtjF8NYkZy0hrdzEK0F7/mywMIVwdS4H/jms1iMcM
4OF6k02HvufPhj2IYCTFCS3Vsg5dVVPQclSS89foWp6CHIaOQA6GUI+vkWtGgqt7
uZiX1AYg6R9Y0YaFHuoa6+W9mG20zs58s8WO69K5wdCA9LvoMu+/e15sddQ6yQhP
0IhOFpWnxzgWSF/6c4EPx9Le9+WOPOK6f4CB8XMt8YZQa8Pf8juaAIj/yEWD3HRF
2ttUpdVvKQpOI5AXKF5BtYx2g83UZAfD0OTtTcYkmCL9Um0T5BtAwIKBshkO1Siv
ZYnSx26F0R1TNTQDABSf6HthczdIytiiY2tKpIB4xN+2rG0I5fXM/cAeqwUljFoo
/5qH5QhNKkxdgURySoN2+2orwtb2CaIRycTwMsN+J5IjeCWiTSWrTuoLnHfymvKO
+cA538qBemF/6DM7k7yWnGlGxAWQFhm/gXRCpn0YHGgw1k50gjvgHAbNCgm+8Wt3
sG0Oip3Dvs/iETkJ2JxPnjnQ4Sl1XyRhTY29sBod5r8w2kkxCEjpmAXnGI6pQK8u
1NNsTRH1s3R71ljoCOlh4tcXvrOe5sy3NvSbFCuaBCmctO2arnPOvzxb2I9OZr/f
FmFsBvLe+597wJaQAFOsawqyZLclimVHn+n8U/u50L0DmdQZvwT2sNmyJW1Gevaw
gGq0IaR4DDDTIp2lXJqzFi1qGf2KLpCPuTMK2sV36XhXlQCcIMAhOWYZInqtAEB9
8ho5wdfRp6ifnH8FLRFcUt87AImV7rx7rGxiewnr5IQ1dERX+q4pleri++0ZZnPZ
Nj9oIzYPa8wMF26HNcYreW2UjY6RySFPYh3SokI7VrX1Jqy7zyq/6Bk7y67bbYvD
tN72CPHHG0JDFhGcf3UYjTUrhBkEhWVk57hJRWHZRLMVetb4thAp9ufp7Ov5eKh3
b/AfMbmqQqvgXpDycYnRJ8ydDyp7WlOOPkx2tSppz0OC2ZBsmvtLDy+kTCd0wV6N
JfFfQhXYGHzfYEAKWPyvo7PEwjysEGxMCJEINkk7Zb0KzaHoziUvvef18jGocMyr
PcWiC5n705P9hPWYzjt1RGE+7VdBj2M3kX6xoRt6TLqHtX/fDI2tSL6+P07+zjSy
BJF76qNIWYQSN30fVAxc8jovAeSqhshB+kGVLGKwHiv7+rHE6s/cLD++J34jsJcH
N97YK6arbKU0Ybbt4msAGdCdy4dJQb7s0baIMvB8MqZGWApRfFFRHyv8MqAe6fY8
o2Lkk2k+zpAwBw4rIspdQWYF07E4BJc6DVUCb1bL/LHBnCEcBnNIbl3S3rXIvXty
mIYPs5knvQSv7qS2pgfeR5fNVEsdfR/3UIdtc677vtQuLCv0uQ7iFN+xoOFXm9+P
cj/Vwod+Wk4q16yOstZLQEd7QV6foKrOFvILIHRQmb0JbRzJT0IOkV1/LQbPh7Ii
hCoRGoSJ9lt4rdY9Nk9tYKllLV75Fx/Xzm46CwRGZ7AvXle8ZhohL58jxuEBlXpM
7scWWmwjPSJppip+yRBufmdFbwTyGWgVRLcRhOVQGxMKhjvl++pi6KGmTsHEGd0y
X57xCI4LD12rppeLeWi1g62g1bq5Cn8hQaRfigodA9cJD+MTA4biWwxo52nXT94w
y+Oj1/59cPjdC4qNovRz3Zm35Z+SjqS+WUMIEo7A7JvQUmAAb+zEPyn2lN4FfpSh
X6B559TtVVBb6TwEHwcuymOt7h0hBNbtQfE5wgc5DEpiCgkfjBsTV6ERbELACOu4
7POe4jPdPs7Jsrf+8CoDmT3V5DvdkI/r0HE3KD6aMwreOUm7+Q9Lmz4AaeiB6jgb
mpS6PJDWMM0kH+p8IaYnsQccxF8AKBV3L/ipd5rdV9o+5UnhgVNbK2re5ugIE03R
BwoQxbiy/8g8CyER7uf+dMYzseAdTYUWX0jKOhFqjJjmJ1S+5Qkmefxgrhh7ZScw
BMNtHRnAdESGl9aESsn8n7f10/6hX+VEjOEdndTJMp6ajPc4UTbT63JCdl74oVL6
B+mLyECJqZ87dfoYiwuujqyXENyTNwwPyxlmkYBirGFVtbn6rwfiakAFBCyujnNj
dzBjYQM1S066ON1J3Rgm+FkcRMx3CZx5bRgRDMgPTgqzntoV9Cj6cLRt4Tw629q6
VnJ1DVV4osrMkJs1D43aSOv6wQhF9KOTIaSxLC2nd4VrWu2Vy5qQ/0o8hzmt1x6n
TRBfPyYXxXVRxruinmq5Jxz3Dgl2zTo2YJntBS46XvJdlSh/wG7Jl4dt7CmPxaBV
UVOSZ4Oej1rgrEBpnHoOAPYzKovCS0ZYaQzHwK4Ugk+QOCHiLDE1W9xrUd1jyygh
ada/f6M+14ojbHef8cJSGlWiWfi96hBMsBTx7ODaWmdOuDKurDB93GHZdKh69JUI
Pmp9Zpn7LPIBRiPO5UBLthWkxscGEig+LOhfF0aWCDXO8qXeb/Pdxk83FltLSPg0
1dpUWHLOOaHT1ZZF5yq2bVd+UaY/pmUri3qdYTumC/B58/ItqEnmE9tPHm9k4r1w
3/zUSivLTZG7Tz74JT0+PfyIPmLbHZQtBrPQn9uMt4EffWO4qoAfzDEhQlDrsRvJ
aU6N7PK8UGDS1RkoOiJawi+Zl8YKeHUhOyhwLGNlJuCsm7WHmqgk6s5O5pYcj9ew
zOs58X1T89NbaZH1EuGHO5yjMgjpguub1/aWDlU3LOC16K+sbDEtL68OoukZ6Sns
FRFADHHPM3ftJYH6E0ikOaPn6UNYT5o8KB0fyHITrmTT+tw+Me4DX9lnwJfb2Rht
TaozD63BTY1LUNtMx7QR3KN/j0nulBPnJOe70s1cdz9zYs04W1756BHIaNsx4HJT
8OrBgFcz1z9+wYjzytiROgREXUll8RCy/yAek6aFRMUJ1W8UQi91SfNi691ZmnGc
1p2PK64SYf4StayKircROOulQsdR49vOerwENn3lk0whRPLj2Pbt6OE/WJXVANss
kwmA6K8B94vemXXgauUyh70+kcQ9IdhG8VBfq3poZMhIozjM/jIiirv5ePpocQMH
4UsVx+mYJ6mtK3JDE5CeKHlcq80aZBp9/rD92lhYQLu7s+wt2QmLPiuUIU6QWjSH
kX5g4uSv2S7v8jNX687u68NxnbyWpI9F1b1VzeZYTwDojtbaiVbX9JNdRoI6zO65
vHwZ+Q1zaSdnbBijyN78NLAhszfiPBB24GYXjVezUWwfIJxXglab3HagOCXwNXNT
4lvwPg7yZ5FwQigVkFVRijtiv9hkQSP3Ql7dbHr8XCYOoR7y8AyQx/HQLWpo1Rsg
APJB5kUjBzk1spLcGWwlPGYiwdEa5/NFsYI3XZuIp+VIXWJ/xO650ZzmPkuafLED
9irK125rZvnsWJafmIkVRssvAfzjqrjXp+14AMZaEmBjemmZ65htdnf1wtbBdd3B
U3IbQgw9wdmYYOdr1YR0O3f1hE/B8eTIJCHWvJFKudmSxaZKxjsvsvmQpcvhVYXE
Lq6+yx0AXENSuivugLFO0hdpxj9hGcJdDzr/QzADzHv/4+9aGdg0MB0J3nUWR7A7
TxIlJoog+OfN4r5i7EUEdMl5Twt/MUJwnCSU2sWvmG4xN+eXDQEgzEoiQ+H2h07p
OYSIPhnkewTbmUPfgFtuwF1nQqoxBqKe9XcgYYtvu8Bz4yYbgjNQ7Cn901/4+kkB
KRQNDkdc1bhsrvylPzIPz+06VLxWss1iIK4D9BY7baPYrrw8Vfs/7hriCZOR2ES3
qrY+8pDi/ASaRunUdhbp1A3MjdGaPIVUT+bpDmZW4KWNswl5MRDySXoSlP5a+l39
pvB2nJRXqhb2skG/b/BF9agJ/yKWEMXXpc+Z2D00WH2QocgrXRJGCYxqHwOhtnXz
ttCJV06IzT4d3MzCScYQV1igY2b1Dmhz8dsIIY1dota6A4EP6yjfMD2SXLgdZ2SL
gDNVmJVP34i7iT5NXknzZNIy2RWH8l9HMVhdevqJ/vYjAkfo6nDI1/3w3pBkAZKp
Q1nsttfZfEs8ogBDokOtt7mIEBIMfrdWi/Xk6NeO8ZD1uShEYEn6R6VvvHo5DQly
2S8OAyNeHMJPcz+RPW9QFRnVaJdMA8L+ztohZuN8YGuV+F1yo9+/7XdBmyCt/TnF
j/yZQOQlxn02qKUknx6AtT/yVQRmTmR7KvkVv836VSiZD+XpJnpKo2eF+cDyI6V+
a9ZIYw+qhhI80bD70hSc+UpiTlI6iKdKhq0gGyPfIWAEzHHMF6OYDAZ8MgFY3/vz
ZHVT7ULmL/wlrxzXFxnhDlrbDsLScfh7tjNr9TxIrNSomtx2mnoqkWGqL6n0eG30
U2ntb3K4wpQm9JvcNHFHMjnTvvK+mUbhynX4O/WuvjoAObq67qRPWqV7mmMQqjwz
BNFuxU3KqMusl0s+8oNP3zVQt2A6bQYUzqs98FLlba0ZnDaUGmSUDJa/ETT5GzpM
T3GqX4b0y3rqRbDcTZ3Jsj6GoH33L3kLBW1yl/0J4fx27w5Ta40T+oRvNP/fqmZ/
jCNEDZew99XyVmikc7dolc3Z0UepqlsSUlD6cR4+5LqQxlxkHewAhe0SqNU8M+DA
3kSW1ccyunGw08EWcZy5QNS8TImvnuiU1JbBWA+f3YWo+du4hY578G9xMCLUdCp1
dpdRr7wLx6v7SEJOlJiJp0ZEI5k+iuPs7H0qPz2T4fBmItKiwyY9xcLSsTx9owp1
/r5/CI1MYz0gZmqoTQ+SYOSvmIkFAiPNBmIKEgABW52pId7jXXouqKiAED9pthEu
bdi3lVPRhHj1UpJ6Xoa9me063j99Jq81jrlNQ6Nl3f/C8cPWYNxRPuv4r0ymASpm
oL9TxsEOiiHUb7rua6GlEC91w69kxj81CX/+SJYPWCel0LMqfj4ECPhdE9S4ZjiQ
HsJnbFR8GC1AzF9jvBV0t1tfDRAFPrhepUhstHt5xwcLBSwDWgOrHvgKmWhosHxm
yPNRBuo8sEriaH6RyCeyH8aQXh9AvdFwSZW9O3gif/3kI/RLQ0VInqplRZPG78C9
2+60ipZLjV1DpFwB+a2Zsvq4uM9ahGPuO8I5NY7gd4T6b2EhhSFLm2+2INc4PlWh
xiHqfV/rPsYkh7l87A6oV1Zz4huf+OtHyPOWvESjjzKCwuD9Yde5fqUNLWoECtJV
C0uPGACZDOeXqr4EW2hNJ7/tFPUgwqyO371hao1CuqdsuOOrxo0gDcf/Omp8SswI
L2M/DfcDWq19rHSJtE/LMOHE/ozV4i5ZrRA0P8F7Rw+xkYfAgpj9NRRYEJWzeZSa
DD64n1NyGxaail5dd3sbo4dCCDPLuUzj1kROcJMReU/3gtC25xhL5SXhZHTZFgn9
BwZ/IP5tOg2/4RP/9XJFvo8+DPWMPDQhOtH9YcOucBpIPMfTI5Ng7qCw62MfaVco
wqMhc79b2NUHBFCxrlyKn32Rd68zrhFeMos+EpKA3wggyEdjkBzWOjbMbgbA5QJI
VPw6DcTK0SiCnh4D8JKj0OQQpUdgCxeMsEP6ZxEKWZklgx7dg4XsKHzyCdjJLX7z
T9qtN5LJjzkq4U+hqlDfpleS4RlaJfPC7sf3sGcSiO8csFCkkySj0PRu84k7mQvi
BUWaYJPX6/z6zX8GnYyHTkmX+6QvB8mDKis4P/t1JH7QB1tBrIsC74pAz1ZLDMOj
fa65DsdPRAlLhbaWrrcBmBFVsB4dN7INoPyOQrc8VOPbEn8pHRVF9gydubfmaRmg
/gr/4p48MUZlrcIoOa92dzQMNjIWj3/Bcs5rcilCd7+bqJW28qOBkuRvnvLtNdRq
DGUpJ77E3JSlKBceppp3VERsetv1GL8yTEl2aU5l9OV2xmWB9B5uxP6x75Dqkycc
UR/BK0JYbWfON+YiAMKoXewZZ4KE26Ony1oKHzA90Pd/YYcRQIAbJCD55dLR7XOD
p8mfFxV+Q/Qz7yNfRIN1E2UaUFMxxkPF4e6Yi0MgL6VfNPCNEx0KCLSSGqIn7qxZ
OlgEPvkGuwxbmTZ9tgqTmm6dm4Nyyk4QimKv92rDOSTMl54lOOklmQCVYyJe7Tru
2QqSwtvJl0nVG+oYnAxXrhOgZ2doF4YLQiczgLRaWZtNtsEX00h2+M8StfwxDI8J
tkR1cUeRDOMv9yAXcwv99CTsHbgYNvm+4SPays8U+1ItHkcW8OPvsRCJzt3DNlOa
pZqWbezF7ty4amTmKVllPaopqHRobQpaPeLZoqhgswDy11O0VvIEv9Y2xTmxeVBW
oxYhXxaHQIJTQhvHJoDr0bqphQq1I8IaAF2lnt9e6MikFCGgLfcwiGLrv72lpHo2
r7rgb/lZOh1fHQFR0rS45aqe/St32079DmcktHVepsOsHhHbCCwO2Hh9MpCpGwV4
/n2ZB4AOhXuKYFIeW8iIfEe2LUyk3tF498yYffDzDdkt8rOvZISPsua/YxegvcUL
vREHuyWcM/mq6t1/a6CdPSVDZ+/cq41W3Xvu4sDnaBH8cqXqKsxjyKFl48DGSocA
YtkKMq6NhdBe4cJ49mIyMxtl4p4xGYkMEIglkBRUj+ShqtwQuIWh4t9Yxp9qHxTB
g4bOnsfxhxsYUljXSPpJt+Q5mIfEPV1CZAcI10aBT4/dF9diXyp2J4JuG9bnkWPJ
d7PoWPwwvoOvd9L4fh3hGvn83Vwit+tzgmXH4sAttuP+3rdZRHodzOwkraeohsid
w+GYIL8n1RMpO/+E5VRkISkUfv0t5+4vQyKMdAgVeSEwHev9w5k5qGRsPF8xCRZZ
cueqJTOqrHNKpEDWlHEevmUFahVpNAtXWiPozIpvYGsK/MwgoJhqsip+SUPv30S1
v0ml6agjmybzaVcK/lBd+bLUYkE8Qx9ZpcbzJItl1Ww1dL1JC07hMplEXqtLdtuG
GXantbba0D1jiTr3v2w058BLYRItb0JImThekFqq12vdIQ3D+GUXGA9zAVl+Ei+P
ExRjAILRkAFQTgK+JXO7npQvn9ruySqdroiVIlQ8azGvHumVhBIMml4pKv/gY/dO
Qe+cNFxLhisJljYwf+7LuUVhBCo54kxs/iN08zWQAeIc+2Ku6pZD4Py6LgsuivWI
kkbyByKsMfk7uJ2kq4dg8ULBasMKiQiS1rBRqY/4UzZS9EtvFw4D3e/54gYuCn/k
e7UZp0CVegnZY3MYi8/gBp/l1Fu6ug5ADdhaj1qpn0yGQlZ3ng7eYIslFiEoIET/
9kxGZctBUJppV2wTVG2tPCUPFPX0+rXAL3vOeNXpmhr6jvXa8zq9/02gucD0Xehm
3k0MCKaDVPVbbc8x/cINeSHhBbcYtw6KVIHw52WfKXQ9wEXAWjROQmxRv7dFrSjk
r343ptAqS0xIRylIRITDV3+6hFeDkJYsyNDeHkz6RehbEM6RrceUxzGaaIRAbz7S
C1QW0HDMhbOZuDtZion6E3BqcvL098tvbJsHc9twIjRIaJcgoka2Fq1VNyXEP+bo
PhgnSih+TPxepZgY6F+f8Aw8U0esK9eTf6Jh0dvu+P1UY7jp5Z/PMfNAq0TLbd6W
WhFWvMfnGBRAN667wpyW04KjklDtVvKetFIczle/CUmxVo9zKLtiFSA0iSV/VlcP
Blo2IkK7uJtf5h2ViziUWJmUcx4MWTRAVZErB4+E6SOF5xv4+s9YVYEpHuNjyC0a
JcyU2qOvhD2MVBr9Yk2TbTro+M1gH/YUIKZhddgc+CvNpFClpDlEX4tHbhWU/gDh
mj4JewG6HAsX5bMEBKmaPz83Cu3LMGelhLHySouastf6sa5DS36kr3SxNTzfrvec
5jmKgHkY4dg6GFjEA0kqI2DlFHGxjOE4CewaPa4NlsZZV8NlywQYCs8VUceD0Qg5
6FnedUBZnykIFNWpquDo1hXa9zwZ6oQu88jz8JLJOOta3FlzEEjUFKh1qKNLP9T8
5X1smkchym9NVBiUTCgsSmkBjkLhrj5QQmAYM4SXJ51BTrx/GDNry+vIGU23OXNm
+w6sRKeKl3jcHFQ5PBQrGwTbdVeebgDT0KakkQ2qbp2upj0IJKAkwJYmj0du8m1l
qtEJPCrDEIXgMDnISDnHd7Jk815Y/gRMgbU2sYVTy6Chva22hryb9fyXN8HvWNsk
97m+bM53YWBRbxOxxk3kZ+oLlvLV4hh+SybRs++7kB1TXv/OV1sYxcXKPwFApEXI
PhT1LElXB6vLGiBY+Sxb5H2Pkn74zsZjMRr6VqIG32aHEj9+gPPxTgTg3Nk5XFec
FmWRcpBUxJ94GTlOGHP+ghJlVnfAVXLu+d+qhWYXi1KAaJkalgvssV3vrr+D3pbk
IPBnP5tRDlUuLxCi82lnjmqINSVn6oltANOLZBHgy7gwgjDk+YzFxypc2K8LGe/W
eRiiBnsTuZjz1/5A1u0eqPkdbrpsxnBl4+ypIglaVnL/B/+oE5qqSs902JaEPBPa
4XBqy/vVNUbSGYXGHfuDZ1Ga99BkGUMVypW8AL17lck+uoYARAgxoV+RQ7/Z73WA
/2rj0Pjcb4wQBsxqf+D9xfZEuo9ocU0KXnW+948L7rTyqpkB96bk99MdVXaKSQlD
lthCMViDdi8MJ7dW0l46ADLX6L1c+41dBNRCBdecrgfXJU65zQAcF7RSIwM/x2ix
RNVCJh+k9M6AP/VLRqvWl54qWdsAumSut0uyxoP0oyClYYaEaWkcRdcSkDNs75xj
J0/FxRwP1vea8TXkUNX21cxdq4w9xRp7vJfPV5S7LBr2XoGd/KGbcH+zmdd5p9la
OTiCqBPpc4Kz0G1MsCpz3oBAHtF03V5vHb5Id/fK3b0UHXXhdAyvuUJGD7KvU06y
ttQB/H39wRj+jLIrwgPvs1qHj7m9TV9K8iL6zTtkvp2+h0STq/00KgojgppkPH9b
z8j/etUQC0ys18JZlPvoFgmYgA43na6qbz2WBCXET9mOXp14PH7qxYWEOt4cezt6
WrorHHAy0HrD3ykC9N2D7MaNnUmkPSHdWzCCMR57SigKMuSHKixDONInKxM4WPCO
Ve3aaUXARi8d/7gZQoCy0wSLuoSjEQImNE2B9XbEfmV+4Sdcuxk7kDGD049sRvS8
QbTk8RBE9uLTwBWVEF0N0LqKV8CFP4LisgKwUcH0sjNM4Ut7XODFzXGPIqn0F893
7VF7w1HwE4TUU+tPwrDHlUzSiMjjkwLIiI4JkI2H//u4lx4RpGvjXPPHSJMGqo3H
DnfJ7R+h2H5wjHrG3Z7KentweKiTDxgDgmVhfQXNbKNbF7+L4LOg17gXDQMHH7AO
9YKQpF3P4lonxBpO4r7xjTqXZy+nUFdoKJX+Sj1a3TAMipZd/RNqRdjNILRkLM1Z
Mft3Dh1ezHAWPdCt4F9nn+SF3/jr0KUqTAILmqizEPtxfR5q6Re3NcHovrvPOplm
JZ4PWAciKx2Dg+uN0kzi9AnSNryxkH/Pz8glMQJvONmZ23j2SpM/teSwmjW6zdEf
7sjQeieeAQKa6LP9RzvHk9YXbF7WLUMWVm9emQtHBPpbCLP67QsC6icnyEK8T27U
Ff9/G2gaCZdM0zIalQZHKVRqaLK43vpNMR9PwuIx8CJ3VE7j67Gile/COTRoBGCJ
Wsmw8UqR6PpNxKjdfEQFqJfQGOHqHwtAo5ohei5+Umwg+OMooBIrgVD4NLofUmXR
HscNsTA5ATBcgkTaacvY9YdkNZTf4GcFtQfYpfZ+I4b6920bZJXWoa4Wc2EemueD
ooPHTNoZThD91y9e+5B2wq2hw2O9CkhZxaYD/iEaObnBB9oy/ACiAjCfkWwbPTN/
nzOOSf8vDKr7Y0lh8iDy5HMv8W/2MToOTrTLYx0rBM+Orpw3i1o5M2xxENrrt4bR
1XnGrtIK3V9LzuAlwEEuQhljWP9Kl7h3gi90j24/lWsDvz6rmIzdrKHYFKrPzKl9
GAJRTW8GJrQkysvIC7F+Apfv1zusV8g1GX5GAwDr5FXMaCRXC7ZLgNjOznoYIjyo
iSTrY5GknPZQqy/VZ49SRyHu77/5KStbx72q7l0MNwdLLftlUtODIdd9/1ejg6+u
k4LuKK/qPAukBcePQo4DpelOO/vNMIoimu82Bru9kh8kdsL9NiGAQN3YG2XEWsU1
BcbidCoDLUHLDTLsGjBINy/uicq75i00E8QkyHnqwk8Eh2M4RQdgR497ME94FGll
ZtVfTrZoE5jxU6+cbGQ7ogUL3uu9MULAN5LHaJqdn4rWPZCFS9mwfYlmE/egyb+c
FfbRNZaCBLKwWCnrybCIGNjADVZsGQwbs8+w3T6GNkAqZi+OCnL6QKLzgsZtD3e0
DNbMyQm0weD3crd8skReEqzg1q2xXAi7TowJKk7a2THYSIAbqxH88fqrp0ZY1cGu
El7dRHRscUqTIieezEgcW2wXc/tXgoCsci+w/oM8ePOGa/ed0woxXhrQffU+a8Hb
fm3yEw7iacdMJcHNiDwEcgpUjWa6pT57I46KgZ+dgc8KnPXHCjpGbhPqt0xbrY8k
lJY9T+X3d55TbiSnDtVdqK2k5tWwOO1WvxXDRM7QHdxvPLNpUd9ZrqOxaEB4zhkF
FUYf6OMaU6a7LUEMTh2Wb8MV8SKTJdcG6vH8iiJCJyElaqUvi2k0vDNq7GiTeCDx
whO0jz/oSgCLv7c6J6WagFag/LDW0GxO/QcbvrXddfjtErGbTpRIFZmnqF8Pjbdh
IVHHXrnLz4YP+WaMXMP93mMQotr75Gu1gHqHfQ9ZSvadjD/A40VdHPgSehU4Etbf
7CvNluXZBMiZA8jGvrw64ukovR+TnZyauzsTAXdMXuX8sAddxcGo6mBY0t93rvOi
ltLmyvT1i3bYNdXRCUgtMIdTijlBl7iTIolGSJA30bKIC3lRlCVUEvCYphprHLOB
yY9gJ1jCC1ISyUWL2eWTngI9mZLfM7XVF19l4zvgWNG0tmdLoXDyEqD4w4Ns5MSe
f0CgdtwbpxOXM9N82sjPHZyF0ixvV0HxUEsZ6FH7mvf+4HWpMdMPCn6T2jhq9htf
ebjR/6iy3v5FSK0/X9OGgBqK69PLjFDcv3p57KJ/14gHQPcw2HFbW9rdT4nbnvsQ
CWUhLkm6Qesk60QgP9It0EoSkYIQdyIK2AwoYYsgybXpdviF0RRU8IX6fkn+Wr7X
ThwMClXWXaaDrzmj4fafmSUt5zVB7lt5VjS13UptVAdvv9uoc91bdkyGUU9PLVuZ
/6mVAS7lHoHLAd5RCj9ewLjrjoqYUjtIjzYn5S35IzziSNtHCIcPg1H5BhlLCqiQ
V+pcxn9zRxZEXyIqfzmC3RLnCR08JBVVxMuLBR+0BFo+wP1IrNdQXFAORz662Azc
3N3XiTLzDvrmlW8k1y31PihomQ84BbxMdeQg5j92xlvOv+hiXzGKHm2LQOM5skXz
lGtGVkI9uVjCe2+yjpnTem7txT/6jFBTuMw0xR3lDLBhrivQk9FzY3pgrnNCMSe2
BCl8wzuREajYPMFWiy8HoGAoGYo0kVy1vtfA5yhHdkYj0OWQpSC2OJpl4bquhbq3
1juNQn+czj1Cg6XKaeOd2eAf9/u6jPvem2CONNGdEP80982PQ3ySzMkTvSAvufg2
e1v9Ub9RoGHeUhLRFs9f4LRIQjFtFvelVKenXxV5AIRmrQmHGFLtjzBqNfHy3gEt
+lMHzQ+2HeT9Jus7OmIgLAeZcCH+BMeRhfW7b+Jc2U1p2mitwrTHyJQd4nk/DLou
ru2k3YnYySQHtzWruKdNsfICmraRj+4D4QvH+ZAV5aj60aaMIiJ0gL8FShMtZzzC
KftAiryw76dZpKtHfrI2TAE0HimdyomCROzPF/zy2sd1JZe6z+PObt8scPa/CXKb
b1P5aUW0dRa557d1mGQmtguJnPR5tWvgqtR0GuWZOAoxLVDbvsWse7foXcFMIVTF
YHfi+cMuQjMJMTnTrKnAf907FEG9kpa6MV9Y40lfRorvOID/XTR6IeGcSEfQ7gWo
1qMnRMlqbpFSju8/7kkrge/NGSWvyA5pxl7eCqpkEhQ3pz8yBoIXr01JPoOJAtdT
NFasxZt1BgpN0kB19x8v5eXF7FrdmSRjjjrJgLRN45NeIcbZf9C7GwUsVMmhfofx
QSp0iDjlOQxEuM4gVU3VJrVz8AU/9BfnmbqV9pSav8y3Z8P3j7rCzuM+evxPTBzO
NIVl+xmHwkrLXHLT/keYm6R+5WlPs2AOIzNlcqA5vARmUU9X0W6rtStK93HdvLVH
7pikwGNj8/C+/pXcAZl1U8fk0wyUIewBrXT8fd14OwMPcSrD3f8BnC2mjtHQMEIG
1A02SMrWxmVw82eO/tPIIIjrjEpLkR5dij2D/cQtFiIHrGk8CF8OewZejqOg42Ye
DvLjdkEtSPAxxXPUY4w/e8EfOWS84PFstxCUNttzdsh6LhVCOZ32GGPidzQrPq+w
dnBJg18DNVGX1o2PYAwLWO5g/R/KuNk+GutDnEVlUjY95F7SgGl6qMwU55yDhVKu
6PEK68hgg3e+yb/Ox3X+vZSdI3a2FUxRKohUkK6e8Yb/+K/vI/E0I096QaYYN0rc
/IscT8HqIyyp5cfvfIlpM0CaRZdEr5oI5mrpbw6dbBO+LDzv4VzFc3+GZS4sJf9z
DZnsURnKnnuthFGxIoEgC0X6L64UNJL7yUPO8ohg/RlJTGeCWMeMnDBVVmfI2fWj
/DI0m/tu/qE5yk4z2YpBn/Lyqa1w+gglppciEfu84hpWo9TQ4MOj+35SiK1Jzvv2
JXHDFYgql3zsHys4LPx5q/uShTz6FLD/Pe4VgnermfiGhltzl5bvLs849k5y7Ztt
rqGau85twmubdje3zwIkiIZiu8FlLkDrv+/hJ7+0QSRvndxFCf6WMLVkIkS145qp
sl7IFK4yzqUTUVh95zuELzB8CkXobNGEYp/J+LM1BXbolfKCbi0VdzBO/nZUsbh7
KQ6rfta/KfaOPPsisB3Kc7QnVGPzSFFH52nNEJ7Ea/sxsVa1H7KMq9eFv/+a2jCn
jgPezhjasghVtSR/JoNQyTFtv6+2vKGm4OiG1OffM39pNfBpzaCYOvbstBudVWNU
ehOPbKBnvBplLtHahpWhgq5Y1UZs9KBMQQkopUicMzZu3Wto00oKliYP0+U1S5k7
j55DhjVSsd9If5sJ3ewYdUh/xigTEtf7rh6GkPN1ANWCJtNtlPZq0AVK79jXOngm
p6lfJQnXmUOYZN2R+tDeQZzplh8LpwgnfYCW+8EW8iEX4oaA0H02WR5DMWoIHw68
75uVcUElzUZYkTGoeAGQHN2KJKqtLgW8/yVi8WRfZiEHbA2gHn1q7E/XEyQtkdFd
5RTWi2L8H43Sp3//BfX9wo5d/JL79dMHm9HHdLK0GXenpJ86DS+DFbc7t6mIW08C
j3sy8v2Ejfh+WuTivMoqCWGtIrHWgoc6c/JPMOPuQ3OAi/GFRtvv8fd9kipBzxs3
U/o0+3Na9BcKRbqn6AZJJME46pPPVcDP8CX9C+1IBh3f8JmnZB4nT6NkUv0Gp8cq
firY7lIcWDV10McqfIOYeDL52IXT2j1XA92vwY1dTeM8PxYAWgy9KD6bIpaB0XvF
Wr6WEOhQS8qTAv+KfUODaCe4/ZBhV2XP9F/s8BNUAIskL6xPl9QzbH2Z04NNQ4BI
RpKY7cFUfu6cm3i8HWdwH1FL1w8aO2K/3xWtieUu/o9mFjbvx0MvCyhkZjameffe
/yalEOdWV+EDF8CD2DfsWD3RKhGD8Xu7Xz7EAHIOipi/c2jFePf4A/XaORQUmWXx
mstYAGPy8VE+/cFDPD1eWsoKnoD7ZBxrnOpByWzt8N3KFE8I6WqGGASa+jHW6kDG
P/Bof7crxR3XhyTpaQlice/N2wZQFoojIGzGpTxsWd2gzpK2HD43YHnf+tIzO3kI
rHLUKI4tbnApnZ+WVRr9/yllWcFKekmXWnnv2Y+V0vfSq/MdSd8on2zL1lr3O0hN
F81BJVVnf6uri36L8yQNzZRH1o18QBrYTRsl2PvnkEBEDL0S2PcpV+Zq608WAXVg
KCDFIgZqWLuwQi9TN45KF7YpGa2eWFPBiBHCvk+OQTjHCuIbyTfen1Ns3Bsh5y0Y
V8fogt0aAUYFZsbJvNtI3TTJI7Ig+WhVSKwcFSP0CAPth7FbHrHmej1Bb8hGNQrr
0KqMfNhpQL3XqcMIQQYB1IBmwAdjVUWENA0zywqcuxBJngsS3ZKOJ3cqgeh3IidY
3HxiYD/fVuxzuOxJT41fUIOIQkg5TF1xuAte0qcedEaoiiWvnaw5JrnF0PzPF2kT
GLJ4m8NbiP7x7hvyRHVWQXUq9oma2jXuNHvwkdjzBKEdJ1jYgMtUBk9u/2yrvyQk
02UJqN25grK3HcmeO1uYrxtl0hI2QvfFUQRQW6D8yFgmvTLKoPPLRW4zpId9nue3
eBq5keTsSBAOvFZj3P3BxrEWRTV8Bv1HRmwdk5XKz9zZKLfIpPaGqpPBECd3Gbs/
qD5jux8Y4mPmBsQqfMGqMHwBXsErnCCAF54dQ8OHzQRHDxBhKFecWlAHvJP5FTPj
6lnOOIEgqFx7OadYHpCC4+okAQ6zzJ9HXWsS3cYTp+czeBhoWckUhy9BOffGqcwi
cXlCTEwxrqp6wjLecb5u7e3ORUKaISQxGvnVVG0vbrfpvIF0B6DFsMxymuI/bAzT
T0dUo9dncKND1uH/A0yh+AQussJ1hnRIw2A+6XgGmZLPD76oD8MFxwQ8gJ8Ns4rA
A13WE++4sj+ZlLIMA5izl//WdjDwifvV5lGTQIl5/hePRQuHRlgD4CQ1dfZPfFl2
8vXjjLmdV9LZvvfkxpzoI+WbLrPNkwD13kNuKKaMtnwLU8YeyQCwrcA4O60Mkmoy
pYnkaNm/A2ouOAb6m5aR+/t1RdX1rPoOrvqBkFWltg9EeGruVM5HTs0QBL0lrnmW
Tt8QaUw37dEIyp4L8q96RUt53yoyNi3H/tU2YwcmG/3JjvXWRFcjPT8niNd8ROsq
jep/eUv0TK7Vr0n1e1s92uKYcjnMiaM5Fb6p/oAxg4itXHVprQWefgQ81nL0D4wK
3x/qcTLbGGL0LSoN9ffR6ykIj6zQkBFAcZOwbaFUzWaJRiHa/hDq4ubRELtTgQeV
5G/mUlb9UfU0ze8lX+PVOKdnAy1t0RoIbtxLDIQYP5YRofZlswQdLCREO1CaQzXA
BXrZmHebeRD+iPLo5wJa09ekGQMS8PUNwXVix/NXpjnAclaO21yWrGK929d2nBz1
qZVnMDuF6K1qMn2ZVF4TliAZxXRkcLX+U/DNdix8DOrwQn066n8fkhxE8wbwzkg7
CBsYVni/bUhLeH8e99ym38TCS43PXvkZO+qHhKsBRMhHsUdfwyZ2xpEFKGxmMUii
HDp8qfH0G2ZSvdXSg3VEBXBXpty9NkxuIvP+sQEbEEpWQvjzkXjoBuis97yxwyzY
qZ/FHdavazLuPGOS9EYEKtRfJR0bniZPEd36vJoRp6gxgqx9Cs/tf9H7pX7RrMac
kZzJO71gSRQvm0q2taJztodUp9KJO9BUIfpcQ6Wmhg1V6TvIzYyr7/obzLXLC+El
jMOqEnH2hbGF4J7W/hcgXa6JWl3f0UOuTkXVEd+GKWlz6lkEARe/GbgWlDLNXECM
SIB/Q9riNCI1rgqL1CChhYxuCsbxU+UfTxyBnr2md0SQlM1s2NxgTPQVckkaBLRe
XjEI9V2ExUPybpFscIV7fvV8ib5ND6hUPL9xxYDKZDrhVg4ZQRHoY03DMtF3p6oX
Dkbx69QiBSVvYZ51d8Gp49PvVj/tG/7tLFOPswg1ZCyUe0UH3B8VV/3wchijT00N
XfrbEBLo1u2EfVNp9npawAXtBV2rFDGjOGUYlk+5ODICdvqY/4pP3XG9hkLFlFfp
9h3ITpYokBE5lOB8uBSu7ehKgP0tqndbJFTzVDTf+UvxJ1IS1ALh9pcri8uVtpZN
O+kwk8vKwBM/bnv2r9+3kMoI5c45b5+R5j30Yipq6+Rm9xaIzw6YYP2NbTJAZjwt
F9wLN0J1a6mVQbtsUaMSVdtKM3i/XED4DxS7ONvlnW+f5UiEnZ3sNmJTSN6/8i9C
POpsSNJC0IgAIYhNvFtdOl/XmH5/rQx/on9X+7f6cgtRSGybicccy5DaIz3FRxDQ
zgfzuqmc+or6lMYtZHdx063ek3RD+HT4tYloLEhgq9N2gY6GvmL6Le/dbiNTO+uX
p0CaC5RpUIrEA2J+We4zlFAuGXLfwA6POTrMNgUZckDfn6rN3HCKXzyZklsbjMoi
4ikWvoATena3X0G7FGFec72/OQqet/MWhYof5KUohksIeKG8P3J/6Uj3rQQen1er
OBqcKQXMv8uqzd/G6L8hSzMJ9PvuSFu24HDVUcLbtDR+hNNegjiR+aOtDX0L067Y
macX/ZllfpRmJF6WyQTKv/lj7tD+/Hn10D7rkUjc0A2pI2SJ+B+hV0PhPDG/EY9W
Un/86orVI8RE7z1bjZpw72rt1Ioq6nz5HZka5XMPrqvzfOrrZPZWnxzFHe9jVQnf
BrJ8+1y/WCD8vbBb/sBEuSXOnDZ6dDX/DU9aS0+aq6h+m4vIlKXTsnOM5A0XSd78
ZA3OHJHGuUjXx6oycAV5T8cNplN9TN7BTFMipCVN06bePS46pPtoYfZyklV5CTPo
GnjQ8HDwEYB3/wv2vR9+2khoGzU4IM+TT+UPPQVAoRQH3iRFhoJSKA2gOWz0Remb
kjbJkXuENhih2SuUYCYEYuSTDBVbud9GvQ83USPgGjDBweb4f3vCaeZbT4Nsy60C
sMvTt5A80mtwSjo0iAAz5fHnBR4MyWtygyprDZ/mvj8G2HBdRLO1QNUFOJ95cCEF
S58n1mXhpRASElOkPkgoVGbv3lrSj8FERME+yYeAiIIE0eLK5MKp4/0EFI314X3a
Q15Lznnal4zsd/4dsV56wcLG9APUwciVeGM1dybIkGIzSarLjmlFqR9uktzjUPVp
VQ5xczSG77mYzivqHRJ4hCKD/+O5Os/8aW6aU8QimyA6gHIpydPv6MipV3/YmHH4
T7YRlKg9b/gVFAYstDwzRd3UuIkzvYsi9dO219OW8HRZXOaGZt+PKFYVNxC4x2GZ
00Au6H3kvEFRX7kOUK8LgGU6irQ8ZVJQfWiT6t85C14OLGzX8MW7a+lMqFQql1yw
1JbfOIYc3/KSQgTs//ltIwRQtKpX5NyUy5WOu03qRCPfpAy7V7twI4PutZk0BeHN
VteBT0utDNfJGqQEFZTxsT8ma1AERqBtUh1qvopkgIxofs85S1g4d3Ge4BDSndeh
M4myOlL9d6iI50sy+d31TJEulc6cwqaMMvdTUM76t3AyR+KvKjtDjUAxYfOXI5TW
fYW07KV3GtK1TkrrHbUBWTGDYaMxjwfIGhyEaFeDxeJ3D6+aEsAI2HuL2IwYlb/c
f06uNcSLJtPAw8l8SpS0vRPpvOpxiNp4JDzh4Mgf/8j1dU0Lsh4hg2ewqzlZxaZ2
aLJEu975pxxTPb5a2oYi4WE/vlAp9/Mnk7xQF55I0Q590CUNQlvhRAalXTxNwVsc
JCmtiWdrWb6m42x0D58YmJNiOz5hEyUPVl3cRcFGzWbMs0ZWd/GcMfBPM/ifZuG6
EAvHkbgVm9FgMVEm5NYCCLOqyS6vKo6XCgiFSvyA+6ATfMcqPsgZKn8KaEi0HyGq
H811EykjnutYvBwAz9Q18c9IiKYIybHKVRiBgJhA+QsvO2CEGcpScsLr0dCdHnsh
X/m9t0zAO5litPhniVf9rHCV6ReAQRp7yihvYyNkPUaWf0Q82tFG+jmrzTNkuLWa
Ud7mPFcOq0KkuOsNm4Wb3weqdCES8DqBwZW7yyZlGV7v1ENZchFWCiKW1RNmJ/Bu
G9z9/kEO1Aqvb6990YxEJjZ8kRMhrK+Q4V9Xc/bYF3styNAx68USJRqSRik0ciuA
9McNM70O8n/l6FQ8X0eO5f9VNIJ/kuGoMyJpfC9DPgARZHZtjjQp5F9GFzGpdIzg
EVAztkC5+FYR1l94r+YKmP+weyutNaI+HuvNbcm50vRFZxviRUQwKwaC6Hkmb40C
RqT3vIGx+NGlVBY74xTjsLXkwaopPeQwLv3fmn7teSV5k1VRICPrlfr4szytvufb
1NK3r29z57wt/FBfXtOh2CIUtTfTqAbA8wgr5bq6AVCJp9V/g5QZa0uCye45uBOM
1eyPOXJE7NOKENgxNdGG3qYlWUTE427cg0b6Km+5asAqnD1dVAS6OpPKJSZJo6ZK
DDcQE/ATD7/9+YnEE9y3GoY+6crfpxPmlH2/dzwTPSWPl2SQzGapGo5Dwg7YMkHw
L8QqG2ezZ1tMUBGr8eL0YSDvMn5Q5TUj2MiM5Gscena+7Wrjcco04HdYVu5uL9L5
xFuqSmWvNqGo3laAc8HPAYc4H1gts5AQFtbElbPOrU4wSmYrLVeUjC86Kk/93c9l
gZfbr20hU4CTf1pDspL9yDZBnLOJqMZJc9zqQvbZnpZznRURHAh5/6HTY56f5tgt
nryTY53Y2NGBEG1PFZk0pQQ4rGg000iCHbF/zARESHmpdsnoQ+qZrh07lTZkA8Ug
Jll4FdsBOMnxp7PSD5obdj0Ue+GOM6vdFqNeYujPoORFtzzWluHcBibgZc/VTb6e
WI5/FtBC2vCvm3Ec+QSzkKfdL7KWkzB7GAnsG7ew0ZI3ucicyuheVC6eOLfPf1/U
IjQof/nzeBA5F+jTw9JzS/PSiNyZewo4Zv4wb+j4g9jH0/85LLOpiwsLw78QQjJ5
+ti5+oQit80aHDxe6rp799hsWS8K3UnLRSIixLwByN9X1jq2sIKgX0huYRpyZXcF
mfYyNWlWodDgMEEMMZcp+6DXXsPYJCZOoWIna0oKFwVqVbzXIqFoJpo24XyfasiX
JHHmOeBPS6HqHqDu+ofeAAwZm6O2rWyUXB2c/i8g83opbC48xabtA4j5yo8il2qj
/bVdEjo1/5cBRhS6uHA3YYJ8hUqsHkIj7wStuF1kWZ9730PB6sbRzE9dazkSO7sI
6ojdBypoes0rA+veVV1d7RGBX2sXAnZJ1maiQmTu+f20G3mVotrUmnb/Ss9JLCpW
7tcxZZO2qR1+k16dX/wg7psSXBZ+IC/+Ahj1NfKYtV5bDoxpf1n4X05k2UZ4tkiy
wL6pBaL7xhmVfp+Xg6FSZ1K/ugzIBOTnrimikIWD2+RycuAj3a7+SjnnMeCnLDP3
4luxV+NzVVxyMlrm013yGbIVesX/9H77lzwBBSXWnLvMOVV94SDQmYBdnfMoecGQ
m3BF/9yrXCpOshkNnC6XLPZIhSkJGN7jdFXyLtmZmmXK318zHU1zdKKC9fiixvIi
mhKkhlS4X0l0DHfQuOweVKt5w52dxw/CUkgrFatn54Z0jijae4PpEUCNVs66Q83F
OqNocFfbz+7yiMErFuegZEMx/hAs95jl/ugBrsQI+KneGyUrhDWUDqt0t183KAL2
IUk98cIA9WIUAaT8gqavQ+Pnct+6CePOMnYrLSdJ4hbmFVwgiyuCsARWE94FdaXq
dSidpFimBE/HLh1zDI45vnNs2gB8zuHd1p49lvWKav54xNBlngPUglNwXnpe55AU
3X8e3yImTu8wluHYedJ16zPcbz2PBVjoAnGJMceupENbX27mbdXJZuI0Tll5i2s2
jY8pGIqNg7/CePmhwv34eblIQsbf9UYQTPoULtnpli6GQIqmuAbrTY925uUXqLff
ECfCl5yzVy6cKIj0Sn8U/IqpjDeFDJscaX/3soFRmkNa9oQR5+l8xzkK9sqZYHqc
Ypxr7043XYPztCZI+dCTkr+dUCYnvW9fwwkFU0lLmsuKtiQSKdk5W48csxAw6Kvh
pjYdl2IjXPa3TzLTqfrSYnnQY5DbYBPJ3fyiHj18CEtqPx9VloAP1YuM4YlHF6OC
1a/4JbVVIZ0CY0L2NUZxBfpGEz1pSihVjR+VzS4VfJmInafQSYhaaAKmz5JhEHRs
SBXg8NjvLxwafvlU7drZezlpI0NcGKawBiLDGZo9yCQbtNNUND+LixCa9Zf7Llkb
RgnWl26cYHFxv4oPWFXuSyHwvxtNHnC8WDnWN8bzJt0fJCuEyn37s/yonOf61jK6
lh6P2bxO/RFhgb0rHSkSZ0/M5vxIRg2loSf/4AtkbraPqVlLjbj/8NHwwFo1Vpc3
VMzDfJMnDmq8mezZ0tmc5Mw7oL8wlAjvdut7sTpJk8kfbHiXPOwU6OmV10nkeQhT
aHqNDbDjiYHwUYrld/9l79LwP8kex+hqA7mx65SVTE1zKeGJ7vesZn9XvkBZGkX2
ylsJIVoRVFuOeDI2c6EqMuUINwUirCqQVSUsOSdwSXCQFwYsKnFFAY2Lza9QDwFx
S82/0tuiuK0oqXfVCl92fOBlozFYjl1TRXepV1lWgINp22b8VOhMvfPJE+ZgkUHS
vBqeisXPoqPLNFtyMjArfXOanLZtRc9FRat+UkzWVw2DG70x8qC5dQyLbVJ+2RYA
/w/otKp+6faVMyoLfWSOIwiaqPz31FiXZqCkzX/OAG2bDxjzkRfnaoXmN30yIOQ5
FmaZtNAZkfRuJOL6V6MXUHMl2wrT01n7TchsWn2wi1Y7OoZvYV/7TmgYpcAf/l9z
b+mcZs/FVNxoYdwxHMbhYYq+rT280uEmMbCYC+QEgUfUe2bNVeuQ8YQvqasjHwTa
srp9dFUtH//LuLNjfy0eMasQo60k+7elPQnhr95Mq2oENvgEXsq4F2FtJnh9Ztt9
OyqgNAwKC2cEFP7YrUZNRe4ShKXy2RUHPkDzZYYe8MMSJVTIHn4QPvC8bb66ypVL
JthX73zfBdNFsZIcTV+uYp8JbRZRnJj7Y3Q/4c4HhUs5Rliy3jsKLP4b8XZMKGPg
xfxuWtK5hnYhpNXogAuFLL4QRa/iLHgALitezJXOSHsQjmaWWFM1Nr1G2DqQPXVZ
hi6bE7LSVKEQ7BM0fimlxLoBbJtL/5PL3jsvt+bkQ2ARMI9X5bd0RBII2LoPp33j
48C9L9tip9tOqhmCCV0nO3wKB/1i2x54DEtElHM0KgEk+w7sENeoEUGIAWeSXiPp
l1jQ19SmsGW6p4wVrSaAF62W6RwMQBQAPa9qG4rpZu0Z5iTU77RoPBMmOxYdqaGG
/fdAZxriGJGNbpOqx7ctka00GCTV13zGi8y+gSLJ+EYlXPRBrxBoXF02/MjwYTfC
i7bsk8WLKLGptDLLk5cYn6eiLmz4mR1qdMbSgzilV6PyrxXUeCIbc0Sh8Iuqw7Cy
jhIvQRBauy4f/AWM3uokud7rJdxXAjmSdK3wlesv9xiam2cpBmavX4rDpoiBN2uU
G5mgdk5d9bBzlmNhGdJtWdiUq4FpvK++fn+ebwhpMNmqLyM3jdgMmSzdLgcU93kj
jQQIi0jKHxuMIdmSdJCMjWD+67CjbPG0pwUqzSAQGx5WCjKZ9pOrajuRo+YC7SL4
4ql6ZY/K6CZ2VzKAeaxgYO0hUcqBesYcNE12sjwBRA0mjqc2997nBVi5pVzlRuTC
lkrhOMfMYkCHeLjM0sHUneCbtKcVQE7mfRxRAJi0fGb6UZB/4tRV21X9rPJrRvWk
irsE3wrjdpbBcQlfH8pwZFlNwYDuMyKMK6QQzfhjWaiAlojJ6GGb6rSQUWbr0UXm
tMZB6Z5PtoY4VPbmjuu17cPJXDMGwhvhifxoHTtqPmotl9ZX+/sjUo+bZPQU3x3w
Q0NlIJicpfAcXqsVN/6R1HxsJ9laqqomT7jtEN7DXDejreoKG9co/QgVbq7jn5An
lx4vKTlfCTdkVsiWjFF45IeLuKWLYI0s0ZeHSfrki5wGcXxrUxsesxn7xvIByJR8
zaSEN1wKBUqK1h+2GSyYV9fLc1mL+36/Wn3RX300pXXq4lU7sHZpzfXhRBiQsaOx
DMk3+JB6nQvyX45qyl00vSbuJSfSPF76NIHA/bIHevOnAR5OAzkcOl30sfWJU77v
drqOJ7FtUogqyHQdDmW+/+XQm9LTLlpeltJB/Q2go+h0F/UcLBvMVkzodo/DsMtj
iACMISwYPDAHrOfLD7W0kVQ6AeLvgCKaH8gD93yDYoDMjYi4KYBMqv2lIymGMis0
WnBlRCBD6PEBnSLoYvbeQsE2UWI/lkhIOWTiO8GoDOG0TACdAkZcxE9Em0mWHqnw
MWFdub91N7vU6d9o/3+E6J1n7BzWuIDdWT+uELBkey9sdycjW/DHsXo8wbjxV5nT
WXVQ6U7kU/tvtgllA1Jj86hMNHtoZQ0/ha/0I55nbrjIf9rYOz7wX97Jb2rHxFg1
dcaXWunKOEwptDphV4odl9snyqQjF+6V1L5FyRA2jXyRPcnq62mR1Ga/BmEaUB6V
/0hP2w9e/sSNSjnfnAM69HWzAclVMb3T9lz3atz1C04n30SeieRKqy/8QzacNv98
JV7TObWJOQcyuW6Kj1TR5MoRVvgnvuhvtRImm3cz2jy5MGUljReEDJcTkayvcn+5
MbgsXjyAOvwldd7hqzLPZAIYOy58qyknA3ZV/sQif4FJzyZQUyOJu09Cz9rvDa4/
vmLyrXC+w0X00s2IAMZwFVxsOdebL5K9PdH5oyPgueLcXWYyIsr+pF/lJdsqnUqI
FyiRW/TNEH8PqyGJ0B+AZL04hWBF+NLpKXhjOK7Y9fzrPATpAsQ4z+JKOB3ktY/0
RfjB4EXLUC3XMud2wxc/6w5vH4z/ySd6kDyLwzy0rUrtq8bGu2aC/kDOjKtwJ/vm
j9+f45RU15RfO5MOXntENqrDU8LBfyrdiV96wVuS/9ia3G8T7tGGnPsb9GcnnIXT
A0SvL2B2iOTtGjHqt+v6UEr50yX2G3DVdmPJCyj9F/8U8MEMCVWdA7f7LIgSRhAN
nf62e9oattZtdTygQ77MECZ64zX5xL3N+XM3bmwhIdupWE+eOR+//FcvZ4qklV+E
gDVl1amCwpD0obYN8RFavfprK3QmqHx+8o8vcMDoOVh2oNjuezyp4QBRb3O9VrlA
lKixzhLqBIkyzm87qBGUvhTSA+0J3BR1+EI4oq00jWOBpyYkzrwwH5HucsA08Zj/
E/Zq/G7kSSjCoD/6ciGYUyWeKXKWndZRuIDQav/ZSko7DthHeqtVZmMdR2Vkaj9g
AoiqgIKPAd8PHbhmCBgySVnB+vUHoC0Q8XmryMPBE8HF360gYp8p45uvM03hsgWs
t831sKvVGk4dTx5we++EBvlzpH/AhlJRsYlMhhy8WJExoFfCGiXnlyCix8Wqk1xd
f5QMdSNtK1ETOcbwV+WVuJ6l71N3+/DgCWwDDrRpZpB9hVgnYc1wpx61+UarsVYi
idLlORfy16fVGc3CQCrq9jey7YB1nYpRsFiU8NkXQunEr08U+apjSMCkYFL0Hr0m
jZnYbpabu5F3tPJSlbQU3Ij+vdjuncsWMGaWUF/OrO6HjZU9FvJglReN8LT/uiOH
363wAqzJmujkuKpFbbE7wetfFydv8Yb9lC9moSELfpYev8riKdwTliCGIwYIJJPD
fBcMcIT+N3e/KlpqpLIAwJLqhBYzeKK0J5TbFaz2vzsyh572CZ318E/steS0gOaw
XXZEWUwFLolwZzqTfl4nhX+z3lS77pj3IANzEuHaIw2hb+lVDgrG/V2gLTEa+OW/
bYDkGTWBab1G7KaFPiHgZrOW6+gMkmxAFsMzY1AqfasZ3WrrYcDOFtroec+tQOfw
a95r5fTxpq7/JJPOTHIX5HMsVgP172gTaEdnHq0GmkNVahB3VI2iId6Jhm5VTL7v
oBudzH957jjYqK5eR2PVQyJRvYkkRjva230/EpVOQLxPONU1+VzhMLg3lPSztnoU
25D9TkCpy7PSFaCBt3gAdoiDl4zS6Vmv3J26qsm0wuzFiTUZpAH93YGlwrFhDRPn
gjQHssVOl7j5lkY88Y0UmMDLPvl9TPKKE55OoOuTjTTPNZSUBnVI8b4h5ikdb11j
HJyjPOAsugJ4Axhrz36rfqZ6L/vo/qTudd8RT1fufy7RCrNXYAbAZYnxNEQFOruW
mcRab55dW5/6eyJl/h5Mi/FIcGhDlh7Ny0KoIRW9DRwwYSYPGoG97aEehoWyqgFi
HtFENEecYS9VSG3Uf2kcF4uv4bofAxJ74NHAUNkhNd7FUYEwXvxH82f5VWU6Zc4/
JXh9X+TCw4U2KeG3jzupM0MVTILzd92Q3mdzw6V3+B9E6MmQIkd51fQMJzimEy03
BoJoCFm0vUSMytUqkmMDJkD42W/Ial1ZRajirmN5TJ606/+dK9OnnO6Ca7FUJqxk
vLbZG2fdWX87jpIjk8kYIqJLn1nnEOTdZcRunlX62xRUyimDF8mADiTrr/Z9gAW2
88FeXMHw6bp0zzEtZWFJeiGyRo90uIt8W+2WIHkRns0W4UieUnVwWiNNq14f9TbN
7Dh/zoTf9jSRu0iFAeQUJE4SHdYhhySLNdV4UPPzT9HknurPRAHGbEJQZVKN6Poq
6ueUbX0cJm22rXR52kl9QJTJL+Lq0l5Ox7EM58mLdd5AfUAwGNJHifBI7eKMsDi3
fMkjzVRZX/NNzSn2bNHIkNWDCUX5mryhzvFosUAF25OEnqVczi4rk6CthuzK1BHf
4VGlH54QFJ2YWP/LUx/YUw5QS5SitqXQK/YFN52KPOsG2l/aZVIhMIElO8Ua5q36
OYEzjaLhxLiqbqEwkgSkwma/0aYeb6T9bmYIv64Xq1iEkVpcOu052iHkDa3gkutF
1SwTLdR+4KL64aRGmw4RqLhqPOVtnkRVPM3ka8cWRtwh3XLWHDOIzVMT7QkuqZkJ
botm8sXzaqiXkjEMCtcAZfcG7jFOd/WLujv750ds4wV8pB1BiYDM+jZc+JvKIeDb
s10ddjOm1eVWanyebheOL8isJQCUoWElYmsb0pOg1sMgCSpYvVI2YeFXNxzxE5Gk
aQCAnxflIagSKIcho8Z66jlQohOf86JoW4w0DYsiRAtnv4vJZHUxdXVrB85Nt5OW
53EVpXbxyaR3l4sEwy7iWUU1TSM7nDyeQJfKxwSvyL8dsySfurcY3cD8s3AGB+hb
y8q2JAsbPRz9T2elDkTOOQ3NpTlMAjrHxtta1EjdZfgyDpIezl/YLz6UvzcNBNy1
xOo+9zFvDqErkhWsGEBrHCGM7BHMCj4bhN1b92Dy3O8d380sPNBk7zhsAQhhEEhm
ZIKMGioc5O4KM9yreDn279yLJ+YkVzP2n2yefWfV7KEIaeSITEf6EfkIWuy+7H/0
cJA/38LUeSZ6yV5pn7+2hZr/rimpqkEhUCbfVCJ+JWi4LDGC/KlqyWqdbkc2Fgjf
tMhKOE3K5/gxaXxv+8VsptCmXhn+XQrNjaTj+hffWd3Jcf1zud+eeBbKVagxN0lz
Zg0g62TBnOAkN/H1Oy6b56GmHpTSqHnnjDP2k0+QRqSdKkSuGUtFfkboc/7r7y5q
QHsiVs2yy475bYqciY4BQtniOsBwDxWViVqwdN29gmmuDV448ztAHTtBXHPIXKX1
d3iqdPeRyqQHMPc4OBGO+kQD4QY441fUZcLHQd6QvyeRIgfrPnTheFwaHuHMYt8K
6eZMJVd1IpLot5Pn+nSl0w+FcKU0s0DrfdKSojjTN/jfPM0zxbKunmieDwUKu4YQ
J+fXveEu9Fkhcqs8SDq80qXwwDb0/eAA8i5Dp1CnxcXPQ4CPkSfER6nIPy7uVQqX
uMRYZ1lt8YMfuS1tuWm2QpvOnl3Juf+RLu6N5CQWl4tUkIfxraIEtpbY1CF9Craj
kHJlION24yvc3R2g+TyapZq6hNxXflZoEoIysbJQFkWGf2V5mhD20Ka5rhQU331D
txLUdQoM4tUqb3HPM7+K+L6qvUcSifNmbFxk75fSpntt7sY3J92R3Wqps4vqIypX
72nO0INEo/5pktwlzc7gAXkB78omdTIaWmYOX2J8Nu/eB8obBUHT7tRYWb9wuBmo
BtvdkfWp8SJGUGKz+t8FfcQ2TUbN2IdQ5SckJeRIt9C7kO//fq48or5ZvBHZCwr2
E6WDugqPcNKH/OWidAs+r6o6IKREZbHWQAQ4j7b8p+bLuRFj8xJdvOU29QikgOui
nU40LdgJgWdpTp6nJ7MbYHEmGs61QqZGAqpUJgy4c4AZF3X2hXFhV3VH4aQbP0Xi
mO1kokZb4XZA1/g9JhAr0FIIPdhXwywbhrzhgsxxf052/NRYVC6jEQQR1YPEnSjo
ah1d+a/utiu+C22S2olG+Iw/B9r2Rf9I4qR/pmL/IS65sU6Vgdd3RpbFFA2r17h0
/x4TciqkntdWltfs+VR2NyZJ43F558DspU5tu6Pvf1HbI+wjF7IDqT7uud5hGta8
w7dNJQQ7JwbqE1/p5T25cboWEtvF0fM343b+RNAD+jgQsfAn2Tq0mNxFk6eYf1gC
CeN13KZaBwXYuf+HmH//quh9/7tpqLgbVbOcQe71jhGwdUfbZ3BKy9+ac7V3QBei
GvAcdispy3WM+IbJr9T7Dv8ZT1QkX+5x2/hiP8fOgdrQew06pJsJ/a6j2gjxEMwP
HWHWp3mwDlRD7600X2ujSgux974nhErunGOJXNc0j7fe7B9i+A43InOQXHcAfGoY
u5KRBX+c9au4Q5EFMDVyhqpKAoOOoicMASs6kHCbn7InqNWkJnV7lKUk7tjFZ9eP
lXHwp8hQMpA0kcfO58q7IsoX56U99BLfoZorYOYFuoad/8pjN1uq9gv4/CTP7m8S
GvNua7FcGX6rlUzgGKp1hqimkei03YgnJ4dyGx9P60SskNfOcElqHsmrHyrsJdmA
ptMMxA1yOtiqN2W8DuGQt9FNAGYVh33GyAtbCZD5Vs7qx5L7p6wulw756kOtyRVX
x5k5Pm2Ih87tGOLpDeXUbhBUClUj0zUrhN4Bgoe3Rtcy2jl/YdI5PAwmNnBSvn8Q
L5DX064riA8QO1QguGu/2GxdRflmeburolyWtDidnteqFvqhvukdD0D1B8u07ZVb
YWJNf/p1VNUtLB4bSIN6GTPKrUqzIqI9SkekWAok+ZmxLT6BE6yQz0Xn4oFBdZ0X
Mak2hMadVhCNJnvaw4ESM0ch5vIkN9kBCuXWu144tiCjKgfZ/wGlS/5d2YlK5Kv6
TsEK8TNTG9YqnyOtdMGuiwuxKHhu5cQlORo5RLXaLZ1tQ2ffE3HiuVWS5JM767TP
veQWiGNGcRFcozfL1I0iiH0qNHMh1E1GRPuTN8MH5TF0VOWIhhTFfPvBVCNT6IPu
S4jxQ8mtPbN3cKIHta+UE+MKxDf96PWyOyNXD7QeECsdP0hXc+sKlWjM0zIdIsbp
V7ObPPGfa7e3zh7LKg+WTWoZeddjHlPBHSBIWUUqSY0ZEfje1G97Ytm5Db/SLlHL
LzQMp8hm8jtBBbmPUgy8WkQE2OwuvTI6NhvHnOOND1dORXnvU9B5Qe3goiLrSMPo
hYFbEp3RxNBrPuPVL2/xm5eEQpniHqoAwwJe9gJ86NXfHSIHttrv5isEfp87iOrj
rXy4mS0SB9DSgFqMheomyBrbZlRg1g8Ph06PU6ByV9OYCgEZGBwtu+ee1WEm9TDf
N1cIaI85aTVAcDFTNnhZAcbHl2QH1nMTW50vsZoxsmMbrYKcmQ4hzb44rpjEZOKr
u3RoWVSyDS+U3/teofjMTP8PzdNVdLHIYt+FNFMuOISueczZipzxFd+JvdL+izo+
ME8yNBmtXouU53YHhwVuZfyZIkW9+FqeHV29kKmgv3T8/s8/b/FkRwpPqDZdBILW
6g3beaiTDKYALTb1lg+/yJB1Ah8WFHe9hxTVddJTPlUx5UBk6rBafVeiyJigwX6p
MTU5YrVz5TCC5o+eOHwjkBq9iu/O4ZZsIvG+pO0UYiDXGqQNmT7DGIpmaJ8aHRjF
RPUw+dZ/v43F1luduLJq+oQP8Skqpwq2jvUlLmHjYncZKcS6NlYsVyFwmPpz5F68
P19JfGk4Whikd3SO97Fn+1svc3MKTCdn/SLJGs28IZ/H+IqWY7PTNSOeTeBgZtcO
DZGejaD/0pNcO4g9BNHlKHsigdYiaHOTL7TxP9KoCpBcWmE64/NoCl3222CVHALw
ht/x3eZodljXxBLP7pnOiYxzCCu5XFbgZf8ez5VzN6KwF8idtmFFTwzt74e1hhx4
v4M8zyl++oWnnA4jElxYgCKs/0fZRPe3Ory8bTbLLV/+kgQnxJHo6LA6X0HFkSNj
ztFkRyxGJlFwCgnEZsYqr9j3pwJ1y3IVDpGSImxzyLzT+O+QVuS9VA92NEZQyg8A
On5lyh+/Xwg8JVpuRuI5RcrRasZxCiAfbjcJ6gR3ahRh8wHiexye+O/yndXoRBjh
yYT0bOQUG6rA73wpV9dOk8S8bz+LTKGG5Qom09iEmuomCwEYvu2uycnJ96kttkii
1uYx0JFBsJJszcKtdzd+0iXvw4P3qtAL/yAaEgjQP29DxxOIbmnw6T6CjDDS1DZ7
+MfxzyTE3l3SJ/uHvZDjWKXqnT0BBgx+yCr30Y2dqcMIf/EYNLXXEOa8qeZHxMHW
CbWpYDDynLYRVlV4n/x2tdjNxiiPcB2vwj8HW91SDZ0VR7JXAKvW79oO3XmABSw1
pVly3kSIuRaF+liZwGsjCleCcsUdYc3/cw30I8hu1Lmkxe7qSQu1pbt6FGXfsAD1
ZGyZLirayADdphANcKEvzBtZl98RsnlCP7ukaMvGL+kpST6gTLfRMttI/a2EH0Af
p3co5NhukFONIk2gPKuGs9R5tbz4Q5lXFH4pJdUkBmmvFvWua6u4nUmzhfkkqZDd
QC3qpW0gKyJdJmP92bWgSfPOE4io16w0oSxyjktjQPiaC8zgkq5jc7G3bRKqcdjk
vnJ2mO56HUpNIVeXBh00UfsFWzGdqKUVhQ9WtumiR9BNAzq0VOIseFS7N4OyqSKg
vQ5tozuKDuD/burQYH0dRGpw90VK3chJ1h56onM97hVY7QJ63Bieopyzg4dzjjex
NS7/S8RvUfmOpxnqCE8IsBtF6rLdRP3V6nqUaneqeVEWIJp3ajKyyDSu5juxOCo7
YHYxC6ldmIgEKGs6XTH0p0pyWMUSRzszNHtnZdqhlrxOrYyu2OcaOXRsj+utS/fx
MA5ryVcjuiQZZIIUPHUFF1h5sQX/bbUbX9mD3fc2PrW5X3e8CXZ771OWC19QYY5+
GCWla5a1JYmEN+sDpKN203/4zYF2nlpOmYwA/50KfHk7QxfuwfB7rnoOTg8BpI+A
UeLf4sB6DAK8d/EQTkObRyNW8f6ohccyrqgHlIlrkbf+Q8HN4QwP0WczvLAJAR6C
PyAg53fF0v4b0hLwhnx1XtveMyidQ+HvxaDuF3SGpKg+FGY4RLKBi8aAkNSnTAZ/
0fu0hSgfxL/CEnWl6cjOWuB66KdfR/Gps/L9fAp56UiX3friiZd/iGRCdXYId+DX
wa629KGkxMicJEVyPCZwEAOEdCARAL7O2P5br6EV2gUfRGJv47Wq31EJzB3wfVaA
kzFdNER5MOPP23/Zs7Aa0Y+YJnt892v+mtLGeRYAGb0+QCPPo/s+21wMT70GF/xp
HqqKfrbE6xTbRfYNqE+9BoRU2DxRrTdmA/EWdAQJhUHwGjHRGtb67Q9zPP9sqVkn
us/v1Rj4mZ3CsCWdMQwBLP47bTYQvGLBnLEow1GIWEaAdrx2/KDi36LIEkqFMc4S
MvfHcYzbXcxNNtDGWev2ROVTAb+xJC55g1lC9IC3tWfeWY74FN0f8n8E6HrSkaIG
56CkQb5G7UYLC/pPHO4JHI1YeSDx8S8pnUvOJ10iqj6Qs7gPSgoAt5Ax7OCjxCum
z0SYkXRlht/V+QN5x4amqYIxGrg5QK73PlOAqrnZI1rhFm66KlAFcPzM7yES9Eej
suZUsYSFurjs7/kXZ9rxJx+n/9aye+B5ggL4g07a7zx8lYGERZKX0D1zpP4iqwcx
0f61f2VXPPQDetOYWJMvSDzZsz69fjyWw+gMdKewG/uyUHPZg9nxxyv2ugZ0VriC
KxsubJc98xsZ7MXbNRzrWy6vJHlUtyS3TqjpVpyMNeGSEYz8/QGCRDbPA5wetrXT
6i4HahRN8Gzu/kJ+G0RtJztk9YfZ2CFV4zoWoBvdbGQAUGOQ/JeonLQ+hn7vs3vk
2l5V8WprWGQfLWV0uiywV9/VOJwafu/oRuJunPzvoPkyGYTbvC1MtSlg2d9zx1L4
OCcm/G4SVSMlGfP4VlfDUy8Buu1H4MMt4nOn6tdIoOJ+dAqMpFRGc8+eOuH5T32U
6Jnq1wKFYfRuzTiAbx5W3ls/BD6Qn5WPe4Xq/SHud85jcjDWwhLDmp0+80Dm3BYc
H9n2+uSLah3hhuAGXyaj/XYtA+4KXzkF3YBP/IFbLtDu+GxN07aB9gTGVYUlcAsM
urUzSoIXgB+8uwtfF9/4bjRoUTHsqyn41ewliby0mBtWYxjSBoRmLX80gb078FoD
7ypcD88vkYqzusCyiFNnHfOHoZHyHtnG1zwbZhRKE8LtT/sBnJweqKN5dZDMfLa7
oFVOgpkzCMY0PwBI4lZGf9uyOc1tiMN1uQ/Uu0JA1mlJQV6NAGDGJrPuPtxY19tI
+bF+7b3lQfJpz63KAZVFUNZj1jWu+alRwB64v7sKVgr3kmBBU6IqG+FNZY5HP/a2
areK9joft4zEPr6neypGAYPuS/DBSB/TvqHrpMGQ4QO70iSdVck32KbWdogZdNCj
99vjHx0vP8uILX/gXxwbaGg0asAjTRUFXWRX8syLeQAqDA2fdMgY/lNCBrK4VkZX
kZmrSl6H92rK6ZEUe36uZ6dOOhGWD1h3cfATkgFH/Mlug/6Kaap3CMNdnAFoBXp8
WL0TAQjJ5LOtoLlKG9kQ9UONIA2nBCBeDnYaRHLuVaoseDqdHRw2anEic9trHRqy
x2mxuJXWiTzGuOneAmlQGIFx0AAlI7OWiwkwzlWq4SWHTjdvietZNHcCi0Rusvsy
W1LCve0sRJNfaNugDR+nHHeFbeJtI5IVylwAOVYwuTV2sxV5/r7wouVQ+AYOrSbr
yNZn9rPyLByMgGyOuF+95dj83+FAWRyCBJ6b70fTjMghgyHdpEi/nISq/zmrQ9qd
WDIzbHWankPyF80A9d9FVktxwfJ2KcFztDdyz0imhENk/CiFDEqoiOwrE0wUNRYU
OefWwSZpf2tzYJWnbVTT5P6iun1CawvsC5UzvqbREV9sI/OBD7o7VbRXYtqWbhpW
UYPcnbuiP/XGmLLL1ldv929JcEb9Zg8rHjAubL60XRwozvKODcyEoLlad/qoN0H9
qOCG/z6VP6cDGiR4pUG7ntPaUQZKnbuxu3X/oVeKNSSUBpwATa0C0YJxAVs21MJM
O3/kWkgrhJbQXyAsIANaFaPF9qQxHa/1b8ol+TjtPYuim5utT802iUeu+czvN7+n
OyBBTkzSlqknV4hmmX3Q6iJSlkfp0/5FksKBZ50rSWUISfMiAWDv5ZHo7hFvrxqI
q0YifwGsi5GkOVj3dRo1fC4cjJoWmIbsh2Ne74XlNpw22Lu8ysMsfkdqfm7eLck4
cWDNEmhlehGzNzOmRUlzfRUx2CSilCCoWpSsSTyJ3vQ7eTufNk1Y389gKtaYIj4G
V60Pck9bXloKzLKa+7zGAT3QcVDYucjX41/KJXi7zMkuEjxQRIOIeuiO34VkWIuC
tb/bS0vKr0v8V4l+3jBR/BiwziFTXaZ2dj0Z9Xk6cDLbCdYNo3VkAq4m/OBLVlok
La9kTXB6dtvyrhrYxpOU5bxNaGV+YqAmXeTc3n8cVPeTWc+eUyPZHyvMQVHTg2OG
EttBvBEOhY6njFE3e9gN0SxW1k+ss7M3egcyaOvq93HodDPOQjq/nV8upMwG/1TJ
AwVYsDV2cadCW34jtmUczp94ndo+zX+6oXr2vjXX/6JwALNkVX2J55dkHAPjkhf8
OFcTpIM3lXiWFQ/Qzp8KYcEUpmCZ8h6ofBljTp+W2nGFUAG9DvDkgW68aZ8ATzrr
vgfqXiSs7VvJxmcg0VP95zo0st7WufQHNjkzIxrYkUiaW1I03U8XHHb2vXsCfs6U
hbPj6qFUfDTFkVtJFJx5PeUcKTUhiWVdo/Vfp1PhnxJvL0jPRh7BcHqDoj+gIET/
Euxc8xjGvF9dLlm9AkpmgSvelweh/kaii/nhKAdeSUJFVaIstmgtTVJGe7JyjqBJ
DB14CSHA8zGixrXCIdhQd7Nh3y5u1YvxFWWkYymkLlQDaIrsVqD8uji0DKtXjxul
f/dVMJMLgYhWsd4kiGV0BsyQOFjCMIModIJLFRFLjVOlucfW/dCriwJhkjteni0u
P5EicbAMBQn2NkiXnjRDZQEOucddJYwmusfKvs9no5UYS2siBZOSKQcVVYD3jVKj
iEbARQWPK41nosqT5W5whY4KpJvag2PPcFJP6u9Qv2mnpgj/nPZZwGQ8tDnX8uEi
SxKfVNXoRXaAnpPFX5gMu9h92iJwobucxrGO3XSgwxo2IJuEEOUUlsSVEOQcR+0P
K5M24t8TAK8fOK8K3hU1eAPNPktejT3kabmSPUx061zN8UkLE0AOf/xpjCgQcTwy
ihzNAt4ySHuqtor743OT/VaYFbLRKViaxd0oSI80X04GMFrX97fQ8Aq85WFt300/
gZdLKTVuw87WkNG7RQ7WGVXoMLOeJ2uQdmJo+DqNMNuJ3NfG3Dk2hoPg8l3ozm+Y
beejs9pani+vMoxlxFD9BEq67czOrytDGoGGwhNt+74xQBLE978L2jKtPjn+y4E3
YoV9A3bTVKakfY3Kuc0TEsp6oxqHZZJz0o8JGcmbQ6L64v9T5RPaM74SfctHbfMl
qQgCXFyYFkVuSFO3u3d3bJm8E7yQByr2OXBemjdzjIwmmG1Lpx8A9WnYGIdIYqU3
lQBWShgqe8EeNiLnJKkQphSZkuLfiHmk8TUoZ5qejiBkXObQGczZ/zOiC/sYA0wh
soVJ2A4EoJ3Jth00mXubu+PyJBTNbHOhaMnsY8hfgNOeX0sc6C7CpZ/zcaM1FHR8
9WEhsorg9/2Ay3WKtwPuE2yPPx908WKcsTqLGLfhoJkBNVjo4cEPGffn53+hBXkL
T/qZlSO7DAAtES76mYlSJqVnGOPxLM1GMO+fhOFoIz2M/t03FapHD75ot+RJvGC0
t9BUK52a6ni2ucBIJTzmOJ9UMDWEPoxNWzYRD45OTDg5u4NcR1sCzmGROYRUyX5u
no+nubU71tBTxqOtuhHiPRVnGrXTN9LfKUMxIjUtgzZ0YgvHydS+cKs0fNOgILN5
UpCEdTZJamN8cRE+BUZqMLTC5n/2eP110jcZn5cOtEh5Scd7joD5yXBqaQhr3kym
IrVA8iTQna0kfuGx+26rfWDsS9TdYmhzwPPNXUMNz6NW+u/FiUbftIgS/W2SRWcQ
m9QaDOdOCVXgddLgyUiOX/6+94b5xd0ZCtSuqDf0VSa6hC3vcF+pUUtiX896FY6K
GFOjVmvLFlQLfbwRpkrc19zgZcacj+RgYbEBzwFOlI92GeCpePTRr898sjmJpWXD
sG7hsophP56coM0zdXDqppEanD0KpAZNcLbXa4b2GeAEq48eWlHAL9hgeXZDdlYd
3CwaGnQUNl6OVYRcxbwT7lT21XC6c/COWTp00ot1UvuZmXkp1ayy19h7j6BOjVYo
Peo/nOYXOab5h9QSc1acsYyB/D2viGVU+d7xgAXbbiIa4pYx4RprbBt2Zs7oTH8a
L7flKvJnzquZfgbsdZ484/dpLz8gVGzRJgtMBPq8VHv/xJbJfLsL1UaDcgDNMtu0
jM3zall7OfxoGByk7QkE7lQhP5iBTT0qDHeZnFXH8SAKfv/PRWd4OcJMMf3zcnf3
otyZQDjAjD42YZbTkakgXR89KmL4IsVi6hmQ6kp+a7/jP3/VLqquahXn880DRc3x
fd0aj14jS+rMXS9Gtj7QRMqIkp4T/VhYJRhbeuzbur5ZVcHGNNRoTBiUavXqR/FN
EGt+vD77qzqFM86TdNK+ylJWtCv6bB4pVy8isr1QA+pQ03SeyyvNVlPbPDkq1Nr5
Emn1t5jC27MIolR4oApsk+zJ7qG0ciCQN9mQOleRlxSHX8Y2VIYLUCWg4VNIpwbL
pDLbE6c9LvyEFhLvKInruLIyIiLgyXNlge86qn90kT+L0cFetfrebsJxVrtW7LzM
6f8T2qYupTWlY1q7zzc5oCg7WvKb/c+eNRxZRQCd1WrILYA4LG0G9RL4b/gGhlaE
HsDx+16higxawdhkYWrSw1oHhbe9N+QSh/+yWz0GOfRZyrSOH3+EnaZZeiLw2OSa
fElUZm/IiKmh3L9m1dRlrBNK2VW9kfCQdK9CWQaKwUUkg5iEiEPlScvVkCqWuOYN
/S/dHSs0dvx1357amC91dKWCU6iyI69YchOmrRGh6yZZIcQPZ8WLmSZRNdoKUIe5
tblXzQMoEhHJ0IHH7pHnBZE/ZfhhWyqjJL3GU201TbRF++TM0T2gsCadCypEAUid
6TYIswWoMsC1L+4ZFWyzd4zhy7KEGKDtIeiKKY1HP7KEf3ZHTpYR4j6AJJN/6Zzo
R+KXW2SS4uKnCh2R8srOC3OXbDvLamf5hR0pAqii1Th565BiE/ODMHEadA84puX8
XHZjp52JZ87XgYfthXoaY9XKT6rSHp/FUNiAYfCTKZCwgwZv8NpZc700M69eqLhE
MZdR5FZ05vMMfNNnNHGgOO1Mw90Jd1ep+zgqalI6JIJvCcaiA0gtwpao9AF59isE
Jl7W7H1Vm4LGwZG6fpJpU3f8wFXK2okjz6HkXoxL+ja8B6w0WPfobYRpr4kQIZqb
soXYPc1oWZc65+ZeRCNlDrg37pz/oPftrCmSBrcCT4EgCEtLx6vQzcsj6swwLJ2Z
UzHe/jSNjNfym2OZ5N0Vh5cdeENhlkI6pRPvI513BrliF7x2J9F4gh3Uyso8DIxi
zn//l1OaK5IyMQHLJ+Mpj8IvcMQfQflVWbnIwVGxPjmRZBet346209+2w4MEDOU+
X+wt1CK+XMGDNi1AA4Espf4VkN8UbDz2cCOMSyBQKPJXLTXviEWBEaxut5JpK1Yp
ARxd9O0kgElKpVAz0SQsC6LjJ0BxzWxiebIyDuIoxAf7jtuFP3Uabtcspksj+c8M
ikz3tABIkGcEVV2aiGUT6EbDA4qIs9ByNZ3+eOPHO4ndJe2tYWXFPVshie1gdnxx
pMe0956gzY7rULVcsnaDMYbRFy6RUubXaL7ou7gtQbkJklbAZvtnhz7AeD5Q9xEz
ej+XkP3VhcgOgYNNrFIyCH26akhVZEizU9v/7grp1aetp4i4cAqoj6T2PMYENUrK
+PQUz0hrQaMaU+RuZlInMWiZC4Uxk9+zDxjoFTCTViCPfR0MD1fKAn7Jsgh4e9ng
vjcJ/9xkp/i1D6s1KcPMG18sKAlVyEv6METSgLzfP2pII73kayBN32qV7u0nrACN
Vna8Fp8p9F2z023iK5A2q3YteYymUnkjpvhFBY6/hRyX8x/3SUgwul5h/TFhYFxx
BVjEbhs8sU9Wci0pEPWNG6P7tFA59NukKr8uTKgWhm3Bj7I/+78fDqvS/bUxrHgH
epsD6ljjrvAeNXUjpolzBeWSM1UdZYqjDK5XW15EVkIDA1wZkpRLVklLtGPhNQnc
2vqLeOxvF2Yal5z8Jz9Jsdhrp9pXJqZ2qKj+RbNQLUfY2LA6XQOfrpKxEqs4sMDa
mkbivkrP2ZgvSoSPqlQHPItLZay9A0KivWOtHpYwgeBBgXPdVODOfjP0OQmoD54M
VtdUTs6l4N+IV5PWv1I9vAhPK/OGLevpmoNDLjjCejNx2jKpj0JRhsUhXnMULwue
24bAwiYkWyFUZQn7muX3gFRuLA5Z0BFuEMDsswTQGbemv9ddxFJx9UXKhldMujFE
STpg3hF/bLRECB5YRukb2x7SHiQPuRWxidrl0jdUGUaH8cgQ6ZRue/x7cACw0qTw
Tza3fuLIh3ne7dpAjTnQEKYZDA22hUAZVju4p6lLZwWe7l36E9HSgyLasb1JETIA
XwRAFDANDp9NRLm42RWGmvfmEoBaZEk0kGDDmEVrzLPgvC2jFiHIVvONBW9Wp1Cd
Pl8Py+PF8c+FP3+LIiBQVSeXpN9SjOtjtbRr3azDnipFT59pZsQ6jG7tXwZzdQi2
/f+yHXAuvoZTul9fHlvLK88CL2fky94fbzWn46dsJ3sQbugnPvvUO3KmsdxHw7nc
tU0WaUvuy4LDOZuKygyiaTMaS7MCneU+VHOTfDUTPwxPQ95MGybuJsf8vmYJfWPM
U4HURUDBKIVYua61sgkeNSQcrCcxf4kGzYn+8THKdX9uwPEDFG4OHrvkuznTH/C0
WXO2SCX4bGUnTTSMHGaZ7PjvkeQLyfGRFIBBHFqGX1zDegA0+kLGCg9mDV4xx2hL
NAkikwGtnm0/P0hO2IXWns/3OWNMOjhYULjIczhXr35pkSw9BdBLo3mqZ4+6hI9x
QIYYcH7VsCGjqqmHj5ScJpo2Ddnjs7VTHv/9l7m+E6AOaZTse+iZZUNADzcAZQhG
oayrdzWqJl0Xe2GLzNuLfhGzYgH4brneKCZIXyH/SM7InZ4ACc9/sn1RLuf9v5ho
0n2gpMRNICv4sHfjWLDWIK3fIlrdodrNbhpJCfnKHIeu4/wYJRhaJ1JS9OWRWiiT
reToFYCqYO40QvyK+g1FnEpmXHfRWHSG6qFjZCIx6ge2sMduxrmvZOl6Kw8eVSIh
ICRir3pgqRIKpwNFM84R2cb4O5/0B3HiANwEuUJXxu4iSaymLLuQ3QTIzgbZdiSD
x0EJyW/LWt38+5J1HmFYZr3f/VCWqhCYZZMWBnKgJT9W4LaOPJF3+zl8PsPenFbj
1jk1NCKjYxr5RZa6CVrJM+a1+1R0GemtP1ADcza4KuxVJpUl8Xxkqco3onbCF9aA
laCv1FKofdXuPLnMLOnb+jJDk7qGEE8v8c3rCahga5FSEnbF2tXai563KDlels7z
MAJ05CeeYL+2kepfve2K3PhlnL0FXX0L+FrnHGEqn+QoHdI4maoS+/aqYFXkYNf7
OZzJ4BO25/zrywiWCbsIxIvGp0yMPvHEi+blSql0vKKSZvcj0/In/OtxYWawjE8h
XbWNUWILQOB7DkjTEnsPSObno3OF++l2aUitSAmzfD43UMuufq/h2h7wZHCaQxkh
wUhyWCfz2/SW6U9ma6U9cI3a02FIkL/X1Gd2eNnOkp39naR/i2//y1OYfHFtTlJM
O5dJjaWmeJNH+0TAzbrpkpSKqt0I9UNBYZj8q0QwstRU1IfTgb7sGJEmzbHkTe+w
jyb6rVOxvMdYms5ZnMLmylbL/WbVwGF0HQurgqHRsBCOwUTlFyhCMXhQGNo3pSwS
sDVtC6eZSjbbX8fIZUsjXVgK0pVszfDDyJZeHepzJ1ddm9om8lBp/tPpLTInBYl4
Ao95nHV54DZtiD/2Hjw2rtGDmUwUCuvCLGj2vOv2BmIUeNPQWRW+E+CC6RNexP4o
yMRH2EsuTasTzU6UM9d4yC2fIjqSWnAgyzvPHTr3B9d1y9gPb6lE2yV0LDCC4yza
h5mGB3gVdf/dsAY+LbCeJy89DG2+ttHO2wxsvIr766elVbuITLMlFxXprInuqrJB
TeQsZAkri/SZlc1eMnrMaiV09yjb2HjRxU/YELKW1aRAj+KkSFdHd76F8XHyvtz1
cjPhXft5aeyEilqkHqyzFRYhJ+Fwj9MOxrkKd3hZR+Dyn04KjKdtVu2LtM1DNFT2
aLnrLPbS4KGKtkgnnQjuy/Fz+8kr0DAtCOoDcyxHXyFmOC8CM3txfFoITaCvjert
kaFoWjGAI++ghNOctT0hyx2Q7snf+MAviVnaJO5YCRmqBVTsoafh/ohouIg7J+qn
cJKjN5gCXEQK9gGnzEH1vBplHo73qRz7TKIdjp+S2lMeaGMP+AnAbQhuHHzrq7Tz
/dD2qNmEQtBNp1wVYgDMfRe1KQeQPT9mln7mp+B4XXI9Otq706XDRwPR/Pe1uB74
U6lxt7SUJFqb0KrmsiIxG046wmgV3d9V5aHlTUdBJ0OIDL0wLwoCqxMgjQAbsMTj
KscrwRAU8GnmmdiQXpu2fxnk5skavIY/Zm6HMghY1omEXPveYHugsGnm0emnWefv
5TN1jsh6Uac0FhWKpQK5lRa0pyAEhG0eMRP+ozwGYHTsY+93YOJVBAZUaLUJAh4J
MVai33aoK8Rc/YRWXIHfKNiKhAh/ycbYuC9NvAWbQjdUbDNWYHWwhL+rHWf87dYB
W5xCQEucPkGpKyMjA7KEmUBIBmFSMpQV27fLlOyVPeqGpzw1t51/KisvzwUnFptN
c4pYb7hNcjtUOqLkUskVrlaKaJ7AOuKWfXHeNC+xQ9g4aDwLF80uNeBfuw7jqM9B
MBrkvE5sSC2jMNX3hX8Q0TQUX4ogmgkJFEydJ5vJdkG1KmHf6ek9YeMKxPIgNpTZ
Wv5ZEX4/H0BXLnVcM+0PbO2idV5fAs0U6Sc8tFpLJyJb9/w8p/fxnIu+z880wBsq
dUzIIzXt6HOUF+uoWoWnFf9PbBnXXjG4sn+Wll8RBwITStmDWTscbR16yeWRBr7M
E01ItkY0THk28NwbsZVwF3GMLvbg/2fCR0LRX58ea8o4Rff1+KS+/Ctzz+sMW0dn
dpAUBUTek7aOMFwh9i5j7utfpgpUQe8+RwU111jPPmGPT22ZEmPgI8350DUZelXU
hjxAXj3VV+0eaZavefqN3U5uV4uMXyb4+InT1UWhJyXgT2rOzBMs8/pJ01eI5680
98TQWaKeGCGPwfZbheed3tG3S0yPit1HULuZKXU3MFaCfznLDKMzixMI/qGQHKa0
xxho1DE1lpi1atKiWTIeKsd6PGhtNMCCpEgEAIzkgN7QXrQ9RNjVz3qdCJrZvV17
HEY6UGIsd3yp85OlV+Qjzsfov0JA7bHAUKHvD5LmSgiGCPu6k7Jl/Z6b5JgdUD97
CLIXSPpNap5DXmIgqNsW65iFjtzWFsDO5xwwRqonXup+HTXkL+cFN57LiYjxJiSM
CQ4T/fE/VAxVS8w+qGzxOhpDbGHR90X+c71EUBPy9JTNCMKjeYo22RswtARPNL79
tjPZzKOPoy9ZM17HUBmvmK3bK7tZhBvFd+NMAqpGzW68AvkJlgiSF5M7pQYQdffW
IcAeN2IxLgUanBSYukGekCDhVj/DVDLEC10jHnKxGFQALUPqFvHnpU8sRT5a+TXP
IrERILNOWjjeUlcF7QZEFZfrlO6AcG5/b0Lgj9D246JlTg5Rr+O1xxhTVkQTlzvE
ZwDCYwtS7hhaZW2M+HmZoiI2zpFBWLCF8tRQEQ3JFXP4KFZQu3k+TsxyMWZWil7m
hE/NFqzh/tZlqFGVhQWSpR55yh7GfC3/lD2SNHZ7dlRzl0Wo4OmojqeZObCOgWVL
jpjrx9XVRUIKtELWOBHr4f22hMqR+oNldzUQUhiwWnACgQEJ8il9zS2x8Y6690Ep
/X7PTmWDRuCII4y7cp03S2egSg22ysyikAxw3gev/bcFe2U0PJwhsswGxjNR+Arv
nTmq9aHa9ac13bnkTFk6jQBD3vkFJKxSEoGvlBezsEXbZ09Sp1jP+Fecb8jh/Dzh
u1D6dMTKiM4On6U5vzvDT0YdsYBcKvSK23AjwBE9C7KsjJgbWdbF4ix6Lf+eVEh9
Yu9AMK//Ckus7wti39ceFsezIjVMJaW0OfNGr1Huma9yQQxLT4jd9B5aXl1gnXAx
4R8HurHnm4FvTMHEJpHbG+y3Ow1KVCG+FdrLRujY9E8bpOt9ZMb2lMa+enuL8Rsr
oi1anUpP+Ccs5lXu9ud40JA+E26uY0ZY1JSiFwy3k+I4bnfNeRwOajfb09A52DbR
G2A3YO/qOGZNyuLYLU+eF+HCfyJwaN9iv7vUgXAEljAdwm0n8Hto/bjkHyfC2bBV
6oJvTa3lUB31iXZNTPBTYRmIo+7sTCZTSG0JJdN4TC+h+zGWj0SYmsbtbPwfi9Rt
Z4ls09KEIgjmewI64stEVSOLgYAbmhZ9bjf4pk/P4YgW0k3/NCoxLTANqlEj4t6W
swaG2fjGrQBxhApIoKpC6ErKkGab3zvvBTqV3Eggj/xdzEUuOLO2A4eTg2NNcfWX
gIu+qRpGqsn/4JdWDAc07kNo4P5mGWocDKMw2v8TRORKUrT/jLHw6s1WqqWElcU5
by8GLTtsCqrbo+goKDAQCrzvgrgfgA1nn8rtgNPx7a/EZ+yzKjddfypTrc6NlsvG
EZlH2cXpylz20mFRS5IOK1WuaMsZMfiGVHWL23DI4mG7RMSPcOenjTAsHOZCQouf
KhYZIT0b2atOowxpyVxL+OwYtGo5vy7d4Im0K/f+XopwhNOvdEVjbiBYEdSygKIi
Bw2BHC4vnBoy5e8Sm+Kg39pV2OvDlHxD8bDz0MAE40Iib369wfU9gMh7iR4wEA3w
ZwTX9ULSuNcep9XORq5CjIkdNphsoQyyDygXnKvPO5jc3zVX5czFoL3qVSyGUase
CM0DXifNRNJxEPmuLddreq1fONyjYpYGFck5cD4VCF1x3noKCr+ws/2V9XjNgelZ
YLqfK8P6B1kMKAO6CzWHQxtYjDUoG9M0wstoMPZxh3Oz/i26hsm7IwkIl41C2zjV
JZKSj0qp1b1bQWjF/oM2tirv3evefUlzbH5HZwczOWFQKtAIkPh8ITHMIBl8BICM
uI22gzZZQRgfS9bzw4hqji0u7v11i9pUGHzfF1jhHAcs2BB8PrF7ua7dk2AHv9s/
g+qDhGbbbb6PVjwXzr4RcyrQcQmgzIn8tBIf9dNKymtgTk2f8GHI1hvI/y4FXuPe
CZu5Ma65gUwpUTrVhjDMttXtNC6uqkARm+MsdGGiMgejv8ss3jO5H9Ry6Rpf+Waf
+1KiHuXl825DllOWvIw1Wob8PUf/sUEqy2j7d3cebrWjHyiCp7CAozQre+jeDv0f
mzpMHUaovmEJcBJy75ewT6BcxtLh8SSMbQ3+FQkDKYfPAEVIQWsQ4IPtckH3ar3U
Xqu1G5uaE3rkgoax8yRbVobtFqd0prn4l+KqJxW5rVkDVdNqqshPwdDpZs4ZGfkR
iaDz6Ma2rtrTdf/OtX5xLu8CapxVNcAcTlWU3HLlJfH6ox7q85IM+20jO7BWFZXR
fY63y39n3nPxqlh2X0+MxRMV4y52bQkCj4+HeJvBmblHn3phSEa2lpEf9VZ/nBxy
8TvZAHSRdbe9ppQjzwXvhwFI3MVs09hc7IuIoxwIqMaMeJ3EkMUPej099SVlJfQ9
Pqz5yFoKUsQWRvohi32JKtKFxBbwNg3pQ8vFZ1Tf9NxytO9xZY9i7sDepLyHwTkX
QkZ5COZ6aixSSyfMF1PRmkVVfTNmtBK924k1ZHxyMvsIl57Uq2YorzkwuUzGyzq1
vg608MkuwZsqfTWC5g6kcDKMjtTuYbnobFgDsXRNxpGzXxQ5c5gZLE4qvkBWV+oH
G6Zsb1E9LToCJVp6cMs5m3gMe5VhUkgrdLeu2Twi6VSnpGpK9+PUzjvahd10Cda4
goFBPgAt7C0gYCccxyXWQYINkg2LS2Ez5fE0fZlXD8M3xrlj7c62bsBkFQlKRoNC
wMFi1XE3gtcV4DkB6we1GDdMD8STxzTwdye4mxf4b9rB+k4Vnl6iBnLTKOmQnEBd
qde+d4Sl6GPvcuXqSaqAASGLPn9rTdub5Uz/edQl1PMa2oxjbUy/9TZjtc90FsLr
yu9QWyOdy/s5tbxohbr1nCIBTItz2KrNcD6QuGlBpLy0ODA5esrSQkMtznjZK+zf
If+dc3jnzrkEvRhHG0PAtsxWoBrNEvHY36rtT7nEh4XfdE7VmMUuIhhCkj6gS7Ic
rnzwKNvMqxek/RXm6nA4CIo1OGWtNa6+YWE5vQUtfAVQYqm0YA+3zc6ujfomd0xy
HFPcjJ2jpGtYEooixf0Bm3kam9oxR83oYF5Uy32xJo1D9ARWOmWh0+og9BuSgQCo
HPUQKxiz1IxVTCIF/5m2oSV1x3vLqp36DTSeEUiLXaqRpbj++lNGXKRnW/Kv6k7W
l9oRXL4spsQVlLvgG/Pzc48rXBpHVrM3CVXWnJJxANTlRAm3GuGr2ZjFtaqN30pc
wlukwhyDcCMqvxytnwQBEuewZ0CvbWBdW8z6Mpzlv2HtARXtkSeREtUiQWdIcpmH
Q8VhXmzGFQSZt50Pv/1IsrFPoAl2bosbdCF7VT7a3SYyW7eGoZRUwSufZA7sJkFN
UCt6BAqYMP1ln86CxP/rP8W1lt5BAM0ihmRsIGpid2dJxszVCPLMM9Hi/3nxEHnY
SQL5V1RMC2UthH2nhU0P409DsG9dOdaG+0dNjPMp0pQtYBSGC/a+SUfiO0OOY1LH
tiQJPIzDY88O+0ZeK0jpVlm+nBAcvgUs5TkOxke6ItZpRlZhhDLOYz1l0hCSLMTN
l8wLB7n/1rJggDgtRS071tr8WzSPVleMl6gi5LtQIhP3DhqcKYBQeA7Q5uQrGNHJ
JYQ+hIZw/A1Xih/47zrSCF3A0agM92sSTLFXy22bnqo3dl5MCg7E56Iu+yppm+qu
9vfRw3nF3rvZFCbkaxda5KtNizENwFibawrs7xWposeZ61QAZS0j11jrW1EIVSXO
iWTTSbItECU7c53iktXktPqdDKQZ4R2KUPaET2Rby6i+jefArsaCRmjCICwQEcv7
+583R/A9V+ghIw2Thz14fGStKq16S3YnEFBU0ViPjMj44e8NCypBHNOOhGxJu8AB
zVLlz1JsQCQQhdDE0DFRvGMXp7q78cpxJ6ddFPz2zpJSJcY3mt5NM0zYv7hSvv19
yFgBg4zILSsfVtRuZSoNoTlCv5XZmmQX6orV8AqCrsq4PtcGFp1uYyPlTrfRAGl8
dC+q8xymfjFPz14NpzCUSx28/SjdZZ8cd6hHcQCEGVYTMWdGS1Qp9HBQnw+Emf2X
oYrRTuNK0XWZpUz9LWCngnvdkwHOgMgDmokB98mr8mC//EGB3S7ksWQJAe1X/2Y4
D2bKk3OyhU9XDQkAuBOTf8QqGOBNV4FpcyJyan2Vs+v4m2iuEi+41BqeAGTHA0YD
KF79cVEj/Zrg/AEqoZvWyUk3hfgD156uXKAJDM4+BIER1r/TQq0KKBqA1QPTPVJg
EnW0jXEhiy1e4wG9FdCzLCDANz1PUTip4j5W1ZKRasxG94ZyOiKbye+33F1/Ywr3
WSMX3YMJljYk10UECoV0nkYnruqKYZhFeSxlMSxcUJi5nubp1t1zb+nG6icuEcyH
K8RAHBNDogAWDMvd5PVFRH5KAk8EhtAP1v1XJ2lwLT5BO9+5dACSMmM3NBZNBA1M
Qhf3TxcWwhTMzZbHslrqOwCkvR9wWS/mx6LYOal9HbdRLG8kH7/yeQbVlYNsZ3aN
LE6WMMi8+VJi92FQZ1usldk8oCJZiwkmzsmaFxoGGtQTnsX74FxjEazaWqY58I+l
uPIRc80tQ6YTb5lm7/uzPGVfRhd8z4VHR/XiwQIqM/e0gcHiQSX5GvaJgJKbqAzS
WUUZWSA/j0fsYxFM6wg5SWwtk1eW7KAoHidICrNc/VzfjqpdzOj/qwJ9Kl247iQW
C5ydJFuCVlole8q1jOVxymeNivXK75Hyee1xMyTWGGAxwr/SoS3wicPwRAYPzU6D
oBhtRbyy4st4eOvwfyystbZbBRZt0JahRWCuaMygqWnCt+mrN6DbcA/Z6DuYxjc3
W+Qvz1grYOHtiXlF1eCMI+VVK/6BbU15hpBCCHgwLYV/Ly4FTtjmeuYb/pI9O+WS
4BVwmYHrlQPGfjBz1Gz6Z0qJn5qdedidYpH+8YBTECSdK7sXCQv6De8WTu0OzJ/0
nrRKmlClo0na8wr7eagyI14vNzIE2kOPmmb0DtDThpg84KgUn/gCiQviEof98ENn
I6pGQ71ndxQ8xslrR22acFEYs2KYVO2PI1d9WF/F0soRrST78m+ZXJHyYWVVBrcc
nv2axRexBTVgsh3NTY9MOwqr6ua3SRij+j+53hKd8+O7VyOwFSO6zRuSB0tw5tmU
ZC0GwdpYLO0P4+sNzwFeerYA1itNGWQTjEjb6ZOaAwSQ6DSjwkWW1kXvYRA87dx1
aLaP+LF8uaV7l0biBYGZnv81+D0Js2YE04bKUTGzLf+vwdJNJ6BpMmd3hrVNUAXi
x8ssXPDxmcaVrm2Pq+i2yj51JmCuxto2TGvUOpH4IvoW96/mf95Ryird7AQbi/gv
zYY7RCM8FVIDr+93kszZqd/pWkIixrGckmUiUMXryZ25LVqqCcdB93WEYi+Y8Bnw
hlJEoYGoG716dbTKjj19gPK67QBl9j6H0WA4vVK9DlCalPq2ZodNT+PlvglqYJka
1UHCokNoqmXerso2gHkeSIjFSgIZhKN72sFhZUk7jbs1dpgH2qzN3AzOV0fsejbo
79mRXmA0VOxR0eerInEvzr2DHNxDSV2T2mv+O6qFPXI8sZ6XvKm4ZNl/p8WFzoXn
EhGUs2wZ/V9pvIAE/DEJV5Lu3u8XIpdCCsTtKDozWoybxafFH6fexM2DFPU91pEK
WmwmjHaLoqX0HuZvBer83fVZ71v3VGpRKD2joihn7/CbOi9UzkchuwHRuF6rsgQ/
0IuxgRrtCIQjMmmLKKolp0wejA7WhwuhPAOMmYMoiN7smPMBYDIIwAQ6famRBTiS
73V6H+dlT+HcjVNlbY1/wS/JQzrNDX75pYx+CHX2EZF6rM/KUhcPg7FV6mkjFP4A
PiqXG0nc/uP/UYaJfGECNcOhvNnD2yFTKcmW5HCxGFu1mYE0cwrETGGzC/MOPjVN
s45msVkA57OBNLQY8SuNlf4gCEWc7Olj25BYqdGYiRH5hZcTVJLtSuR5aOdk0STO
RcR3H4VugVk6B5eqKU6YjPahhkCCClQ2tNmaA448JDmyZC3KmrF8fA3RG3pkTaav
AwNt4nQiSHcfrEYOiZ1ozZbuBpDAW+hv3JlKkw5XM1Zl0EOdqIR5yWBjnIEQUVbM
IKJza0IDbjwQJ7scjqyyi+U8aJ0Ho0vhvJFBWTDN0l6EIxR5Y5qFjuXcKX6okcvB
WdmNQYFF1co/r7THAl8s3HKkyQMBhmWRsDqsOPB5JBwGOQthNSj1/ZEjEFnuvZ9G
8ApDyMORkAglwqPkdD8r7tJCzoStJmqqR243B3AOrlfMZkc+kmk/bVfiKxsHv7v4
R0Q6Im+gu+qRPFPBjCTKEXj8pJDnZh2BQRkMlRSe8LFR+kdyacNnfGqS0rKRY3pi
A60qWV2jOI9/MfMXueuok4Dwidkl0Ifn23Mc3oxMn8HmqUKcqNrr2vMTO76s7ujh
d27Pqg0P4XeP1fE9VIHd3ubshTCU/5ZD/AWZg/qn5JIENRhEMtLzbhc6BTqz6K/n
FWHVepnRiPfKFMK2eeTiJGJ3clP9eLGhFJe++22kd7/dK/o8jorfh2DKdQQIQmq0
JlzsvcXvC/DxXfUtBP+sJex9htq2KsA2nXJNdzX6bbKgj9aTPpD3vMBA4kyZsCIL
vG24T2baCOyvR8KyZ5OIk22SFOQu7RQ6eoA1X2b+ORbX5E21Aui0QiSf0gBjkeV3
R5T/mEV7VewJoP5YD7KBPdTjJHGXh5W/yHuz1XnQNibxhpcHZ4bxMU2kt+zpZ8tm
8yvTfG9VIfqD6okUC9RlNrVAXbZL54uSSL6vW2X4Cz9cLWW3yMcUqynzmbrQ5yk6
EoYU7XE6Ck4Zz8rucUMGptlRjWsA6FQJprEByYKUF+GX1W94djydVvi/vVtxxYmo
Zwo1wZf76USuC2j8vRWI4/pwX4reO+Pe0JrWuZtxt/o62+G7dN0dH8EYQZuMzBNm
4L7iBKXpg4cWm/nWDkE0Vr8WAZOMTw3rnNx6VjvURv0eod38tFoLY/USEBVovcS+
LHoK/Cyg3Sui3eCiHRguLgAkg5upo8RG1iPzrSOjNAzpr4ZFv7lRX3PHwTG+iF2e
HUF8fcC/+46pBm7BN+SqgQ8DLaXaCCg1YUvjWp5mOrVsx0FSESLO7hEDiCgyP0ul
T9vcsUQzkjX07o3MEQDsMaG6y/qUyEsqHqx0NhqqW1AebwoUVjpFcTikc+sSn6r0
pEdf4lL1+YV3PuUck4ouEw0tGb29VJCjMXiszEbHOk2UFF2QtRTNXTuQoNVINQng
beIhJvsW1YoritianQerp0gR+ih57/9lCaASsfyACIMQjp44dhBfk5a67qea8qe6
7jmfroJkT8Xon8xKGv51UKliM2ChCdALy5CSp8X8XOZuZMx1/oSiAk5qWSzeRQdj
zYfePNWV59dKpakImCGrk0OJszr7vIeJz/7ykiDKiXAZmRe5e2RVMz/nTH/iIjAx
H/Luoute35qDJp0Zy4q/xNw+L+I8qcJBMK5jmI9CxYiG9OiwiwjGZVyoOd3az4+w
uODI4UGBf4tYSpPEPuBEBzfkPrj2wXStGadHwmbtqHlEH3Ylj94O+4cN2prf7IZ/
NTvGHECp2/UAN9sycRxISyLwU7GuFmhjPKXTiXRbMEpFYPeS/9xT5LNO+gk1+XJ7
3TVX3nw8Vryd1/DYo2ZqGeuMnN00rJm2TtjcuR/IbjzZuynL9p4l1lpoIZZEDX9U
xI+HrMXODZMDAQzi+nJIteVMGhK5tEQhLnR35Wbx3NRihVvS74cTBlXnnF4adLja
TD+FFlyxDPvSHJBD10XUDuYw2d3M2a+BomLXviUuLfK3FZZzQH3jnOLl6J08rdMn
mbtS0OXGGCEKo/B4DMchilCBAjjkznS9q1ZAx1sAiToHVY26V33ia9q4oV/7FVX5
o4tEzu2jjScFzUfGaMRHFOZ4EWeZ//Us36pEYPl/NGEhAndCeY1ofIAwNhmN0y0l
7nZCMlJ/4ppGfNVTBAwTLSvJ40FRljz8V9QKA7oqJCCeJRYHn/KeC920A0tBnst4
zxYAUHE/NvA5e6rPyU66ZAOORJGb+nkmMOt7LSfHvSZQudFFnekWyT6IdAlvhvws
5fMnudUYNpLw+aEjuhVAxp/GXNZ8BBZ2jymkKTeFqxpENecsEWDyeqEvuVO21doZ
MuFimo7lqKPYs2ch0sPp6mKUfZTv8/gGX0WR1FJIJwhX9BEbMe49oa0Y4/DHolkt
W1TWQpfxHCB8BwSRiBk8YQArATUwp4xDwkWKBMKiWLLC+47bNYtjXE43sjDjNjMT
A0hF/vi6sEC+p0g/VY/8vDITgamA4W3pnJsMwv8PfkUEUN37DnpSVOrUgWGIpWgH
7NWuqu6d46q3ZQgd0cso8oYr5R2+tjpHcD9tszckhiyERGNKfqdS6ZQlDuwViFW2
zl8ySQG+ut/0H5ArAbLHSZgU784bWnnvpVvQUmyAqBw5v0sAtnFOkDViuXbNNCOm
vxw/qXv2FxGS9TzkShckbFQZaG1Tb3BmN/lGk0N44jP+66uRTO/nABnIdS+UBPhq
UcUMhxKloXnRJnIZ1heJw5XBVATRnsF6KgebF6j1fk1bBQyD9GUXb9EjdLqjCb5L
o2oSv5zr/lT7OgqGgOuVez6JyU6S6CkO+lFnSPZHBYnjIA8knfc4OcWkz65wSXA6
PXwnwhXZSKYyEM4xEb16LVjmt/gSuX4b48SHW5n4vucd20QyUKudBC+0gKGlnw0f
wI1TJUuPhpZXq5QGUKW2W2mzypohtaQAb5po/XJlqb+bTZszIVOS6P+3la2Wt8A0
Y7YBfSCUJzX9Y/DAi5XDSykevsc94jaK0N9Cy/tF32aKkIv7YCXQcWvifZ3JZHjo
+CqVcbrk6qvrwCYeDv7/PSw7x61HNSYLy6aNhNB4Xwn33VkMcIzna9AndGbkyWbl
UkQhz/1DinixolvsWHiyskUvJ6HZi+EIsaPq9akuAUV7OozowCSKwCgo/ZCtUaKz
Xp9E4HoDS8hWo3qvI6C0caTfwNfyNsLdhOy0KIskDsP818VFpr3ijCJT8DyAhE8j
mhVzOhpGUJT0E/u6+oEApr8NwSzSEIfXsNu1zDi97ilbIBGlVhyz+5zM596gkBS9
kLVmvWq1oumcaJdkC7OtBJlXtuTWJ5uobaur6BGsbEL7IVF8V5g7v8EVWej2/YEx
bQQMfK0fWz/PzBO96S8OAQuAv4Uybip6KeKFnPMgV+v2j+gBSkn+jy+85BPRHMNw
bWQ0xhFU4lYigqrWzYBjfJyHa4FXu3mKDcJLzgLEg9hHJQlddBdw/iAHX2mUrtAx
eGiwrhLC739LUASI1nTIpi9sJvTn8ikqmBNvHrk1XtTTxhcBsgD2ec9fDVqKk0z2
zrONtlwYpB4JC0a+8HvSJ/ERL2fb6gSKL5pkH/gYgUXVC1dzBbhldO/KHj02nNpv
+L+cQX6QwCyVhfvFPfWrw7igPxeKYa2Hp+ANTXriKyTigP4gvkcMsk+epXj6kcYn
z5bIzzRhFko5EY4Vi0STh6UZR2IopF+xyYxXTXVLoqy8YCimKDD62V9b2HbluBUf
9nYIV/r1AcFD7BeiYwKOMqbq26bAGDFsw43uIqT5402I6Hp0Wu/qavNjTUx+m9e2
wIl9MlA5N8vpjMPcBEsRlTMSohT+vtEk0h/t0kKNpVz1qZZ9nmVpeV6KH6x05jbb
N7+B6xKymXwJ3ZvgQNfJqfsyNix6V/midzuBPHC2JWJFNvFNX6KSukX/Y/j9X4w6
SF2AmEI97SZHmEFgi65En5xVTPgNlTgANkP244BOr4UgpqvpSWoLcK3s7JFmVLV3
GYTeQ89EJuKx3VrpOGLGaTF9rEPT6CTAgwtV7Cr7nCRktVJ7oE2Trpf40M0qTsg5
0aLGYFotCAsDiBT2HK9716bsIQgU9Zxd/qQM/sfR2MumWu8vxAfjH/UCtw6Hsrtn
sHv4pD/Xaf91mViL3Ur5INJ7WMgu07QobgcxyMFFnK6PyNKj5ogYz+P+b8zTXJ2b
IiwB+eXPxut8x0XsoX3aY1lq4n3LJFN93mqauesnEJj/rkwAcWlvn32yQwGNncMi
svZP5HKKzm7S+sNfbQfALFcngoG4srV6/jqCg72tCuypEfv0b+3yCVCGV5g8DWBv
fMw3ZMuMVd5uk1U5yeh8p8AGCMsYMYx7C5Okmoa07EpMZ3cQmJqlI6+hnzNvwe/n
MKgl9gIaHWywgs7GO5NpyB1f/7gW97NXiObnEvoGl4e1cfUTXbbdLOh7/XOaJXoJ
ZVjXtwYQtE9ylG2HonsBLve92SGl7zsTebs8Whay56d04D+a+gtHdr/MLM5pPAIF
m0hKyt4pCgqxuTNn9VKzPfNGtI4oZH8ls4P1VlbOC5UtEkiYZncehGhDPhWc6jUf
WQQBhvfsh2PpD5Cfvkc+ODtqxOT9QpRCxtyxYZzatgIK69vbHR9aHY/kfj3bpPyw
W9yBxOFQYpas2H8Q3Wtre62LNRQFDUiIvwCPXfiYT7KrYqmTtAf/hdlQWd7k5hya
dHJ9R5zba2tAMBX7ICVSOXS5HDmei9oh9XG07W0czQ8giKHfBBUYuZhiXsiM4ovM
qEPt+5XBZ0mcD6R1hPML6QN0xLEPDdkvzpz1thODzCAslL5Tg/FadfHDnpYmkcmo
AhYA0iRJOn1aFnMC+5oHo/PHUAWKRgoyoRRqlC1U4ARJWfklntGJtZQ+WQHas7h6
EOAhBCq1kC4PhjY90zakIpzjjxrs/uq/7juAXz30yVAGqJ4dCDxuzRxZ7vuHr/m0
+A4mRzTzOmZlIomIcfqz/kZOfjtJ2dHmVYD6H3r1TFM9bAbht6kIHIl/N6gjFXMy
CnvTHEA8Hi8yIe1i+A5yBVyC+8bYcb9+6rjrEkbZv/v6IFabwAN9Tl4rFIjqleLq
RmYf9hJK+L0DsjLEJi8kiZBk6ByeThgYASsdxnZJ1uNIxjiJZSGD4QCb7vPFHC8N
j7lFLzEsOSYIICk7oM/ZjPCV3Lsq3zuMOq5KcyEhdyIghf0TjreHsUONR1zO3Kt6
6LpcG4ieQ61uTAG7LqvbJi2Mx0zGVmc1agLb4uhxhPiqxFFrsMuRut2VQLEXHuBk
0HOpEpBzbdG/1DPW4qkLvUp7yJSCSctJLjACoFHXJOd5ImkWYMWAZ7FyIBbjoX3w
9y7+99yg2wOsKvO7blJdeGpElGQ/7qWF1nehO/txfI53oHcOat6xq8Aif9vfX1QJ
MfU1zoLQiTbQqW0BjXn8ATtcW0YTgWah+1v7lwWnamM+umB3bDrX1yD0mUPc/Dp4
P0En1E4z8zznZHZTXXSL6mdQYC0vtfdBGJUkV5Kco6ABJ5vsChm8dWAqEVucvNPp
HL040PZuFlGZaesWaQnCKcd9niVwAmBxuy0H1YyTyQ2ePLjY7Dwk+5nAfXEECZx3
yzfBA3Ek+vb7R2+9PATK6FgPEQksdQl0kV4b5S5OogJhzn3TUHWn8WHbvhLRhYJB
dj7NMS3l+mBMtZESRL6TT4Crc6P2pgcGS2bH9BF1ZR3H+Lk87vftVR5E92iP0Vht
2BT7ODEy9aP2D6NRJ0cp4QhUCYOSAGLNRxaSWF/OlJEabJgGAcPUPNu99liRCk45
7TViBnqXT3+VTcFIysovQIf9VwOMMsM5ZlfLezzTLubDmiyhleSav9Oz5er2PMGk
NhpY6ylZjNhDe+XFuWpl8aTBIR5gmMwk98RlGVoilukwWvVcra/e+EeXZvm2gXDn
4dtRvCSbwQVz3dQNNwrnZh2S6yN6mCAoznefbRXuRO/F73gh/T2ZGv0ki0etkRHy
XvXGL8tVJR7cPtU77Il/K5fzP7OMmN7aauSJXKEo8DCyytjyL15NUfrJbf3fjuk8
dPCXDgbAh95dbfZicbHqB5IMxlFzZgWD9DG9oI+Ng6tysd12by/Qa0iTTsKYP4z2
re++I0kjK40jdjeopBXao//9UAiVtcz7R+ynmNKYnG2VG/R5zgjQzFHnpQwQZ2Wj
LXS38F19OPzDTmVU7n6isZIGSiexfPPWWWGd8BvbEPViPNp0GZ1udUAqElHNDXJJ
Nh1LV6m2dKXr0BlX2YWMxbAWTfbfOrbE3SHLWRtt5j5auUBBtji95K0d+/1874Gq
gdxolznaP5X8LF0tL22fSsSyRycuY55UkSwzYpy7DS/Kozjt7wkmzJ/gUGFbf5XS
Fb3SjLsN+ZvSGnl8E3EFX6PSZKmsJ2JnKhY0ZnuSpfg7a2YkWYpnnEQiykPYAQid
iFMze6rnNgIsbWjq3z/9H2DC18jDk56AXfsdCzJVOE8aNjalt62P1ZEV0yQkMUbi
zDD4/w+B5QEd8hQTduMzePZthjbxyyR9AGMYhV3FIvhT79ey+qxndLLGKlfxJu4b
FUM/qg+E8kdfUdaaLW99EoSJIBDg8TEgH8sTDT/FsGH0YLDd+AxgHPeH0IzByDnk
vsd3Ml30jM+TX9kFUxNbuzR9YGVoTVRyROzzb2oiU2pCTBe0VpnnOEc5MqlyuQy/
g5aN4ln6d00OuH5J/QwsveeqFjCzQvKGlH2zD4MQR0K7V35tmo14J23/yrbHG+eO
ZFiCelM2vfH4otPEQst4VRDdvUuKJm+8QdfIsi7vdRfbkdbuyLR1y01MxtjzqThy
CCUhuew5YSp40IpeHd6tGLoH1pnk2Jxnsh+ha7RWHkpZo9y4b5z0BhOwAtgvZAcv
cSOR4vcAsu9eAiFRektyFx0vDl8pO9vlAa3t3eGfuoLHrVeMHYPn2B5hB0pububd
we4lDep0PH2jV1fxBrXV5t5+LT2UV/HOyk1ynL6gxyEiB1gphLXO0s91CPaKqG7K
vO3Fk+4fBYFwtlrCWjPFtb8b3ImYjkCzii7kCKIGeB8pdICMbT3gzYpbuZuahx3J
P3tk5fxE7JlXcZlwPU/MMa7Fkz8HG/ju/hzi1sFOOOPN3ZoQx9QgUCVEfJHp9d7k
pf7dSlWFXEqWaB0eMwJQ50dxke+PAgzMdd0qsmjgabSCcD2eyQptsClDfM5VpKso
SGNP5iM6yqcwbzb+1mP237rDiJa9lSD33ZpE8Tl6ewpo0+j8r+TQC46RHvw7VZHM
sc5rvwCRssavKca3SyjHeRTY5rbAbWEeQ6cbKr+2VCJXGsl4R0lNIScdsVoJYZvC
yXB6U1WUL96SF5YNKOQaUpXM/brz8mmUpleU0VCf3HkQYtuLRikhd+x7drvvEEHv
1glXVA4Wx3zzR6Z7b5qX4IaFOFqG69JWS24g/z1IilEPBztPyAGaz6dVBDtBeJ6D
qdsb50933FoWJTfOYMWLvuA5F08y3OsI+SpGCdUbfCl1v3HNukSINBG0d7VIa+xM
QwV+lgMzKx9/Osyv1CC2/Ikar/BeVJmiNbhU/krvhTuFYxRgvl8AzDJOQ8Fz8t96
ciR0SXGtHsogs5bTe2hpsZ6F9vDfSNNn618ZRB9/iaZgQAFKNNkyYp0AmrGHpoIF
3OV9xrL9F7rf6yoboCRTNB78HxqzuKszQo+HY85BgPUFPo0IEtotg0q+7IZ4V5Ys
D6Sk/uE4vqRxAsN2vd0lxw57GMvZDL0SzH469EJLjDayMwvlMgjItSJi/BBdzbyg
mH7IAg9gcjWPXIQGVtdUnCgo+7U1S2zCUE8TkukIQAuvqGhuKLG7dl8+9avhN2d7
OHCHpBsL4iX0wuPfm2NVr5mxcxjxU5pZHBFTp/OA/Nyvk+VHX9uuRW9cWvzf5vrU
IiOCITGwseV3C5ggug58U4FMU4BTsH8bGkAaU0u44riBL+HacI0oh5gJc1//IX5T
CP3MxQQCkTfI3tC+dEgV4gPb8SOMTaDXNQ/8fa6Yx9FKJQT/aPTmgv3ANw0KPxgH
X33RJ4kZ3ZF5O9evrkER5ywp7NvBpZQ48P2OUeFsmbu2O7bL4Bk1iyZ/c7jFb+FW
s98ONzW2YbTMI6bDAk7c337exQ0vcwitUZ8Pjb0rbJn4A+/Rsocpy0xR+d+S1f5s
wf0IPm1TwefGOqWl3kF4a9j7AdprEGs61rhcrNwo5lLmoNEVQu9bmMrasHhfRnc7
O/11G85PPwhIYgAmqv9EglFFTVaw9KuLK9IPT/jab3BoclkP7fYT2J90yaC8uV2h
1uaSqNqt8iLRJrRa812mw46/hAZFiJIxJRSwqTmL6MyU+Q/iyrWsDKAwHgVFnxL7
JaYY+XxI18+uqIkPhwSdpDnCxDFdzvc4Ffo3Cyrl+5M0itof8VZ6rsTeeXgsrz+X
mvJBHWN+01IZK4sst2HPSX6nbCijgYSVtIaMrmEIK26jSmpb4RwmcgiS3D2tHL7W
S4xHmuCpxdFu2y0PB4+6G3+FH7ledMSfPK0R5ow+ulJy6MBR8FG8DcB9rOTHuYJV
Zh7B8q7Nw2Cj69PC6iElpydqEWFEn3DDk4a4IVW68Q/LCyj5Jh1o2V+5+Qfzcm1A
g75vvTV6ten2UQEAuXevZN7Vj1E3daKqdzBwITRBtEz7TCr7mXVUUs33vxDmi31O
tQllp3rqo3+5yi3IZG7X8PtsGr5EtC23ZhuEyFclSGWuGbxLebPYKmCVKM7zTdq4
oU9iM5ytFe5v1vbsQwIg/54aF4joqd67aOLd31LudKIgpSjFpkPNTc0NVJXfqSCh
wzTbQ77BATedfVkrM1ZDcwZk6ncUcsGpe8C2aoVn4aDjz+DCfzJezxTylTLjJzYJ
KgElsxydqxrXDepabUfkEKmHeo0M+bFLviL2KzKgSPXe3JJ652r2AnG0OSc7riX4
1PaaxjWGcKsnY8krXHiVinY5wWx69r82eNQNhoUR/iKgenN2IW06tlPc/QLjf8xV
N9XIhcPDQpQAx9UoB4+irdslqVnA8LAwDTHtYHPxUbrb3FITzb8oUNQelI/iMt3n
63bSLxKWbCYUi7m6e6s5VvXEga1qhv3C5D4YeD9LJNFI5aBh9g074vNAiWhcYROD
NQxp7G0GizvrayLMchjLuZNJhhCcSewgmVwAEk7P/asGDT8Lab/d8BA2E3jH12Kl
dFHnfPE3MGPb086GmgOkYMmga0ApJyQSQ/pEatZUIlhuj7W5oIZ+C66SHleOggnX
LY6Lr1ublqAjALNA4gJJhp3uOqtazmSQNjjqZvAFwROJ3V2L4ygObmW/duSiimmu
aYbe03yK4z9z6UxcOALhViFc58EhcBdaq4NhAdY1WlqXMXb1KXUF3e1TsBSplekn
Po9L7fuKtm/tPmFKBSrvMBIWfn38AC4m/sGPxtOmrYk0L/gzk6TPBDG1m16m2Haz
lMSX4/vsEnNu9c1J6X1oZ3X8759UZOoi/L3hTXzKYsN94GVq0CDCI7xvBAiyWHAe
B6lZHc3Vh5K+tjXOALXZyvhAO7O04oiW/vNMAgTLXD8l21QX4XEY+NLnhadBmO+6
BNCiQejNNrMEaXqtz88tgnfSgoOEWHef0+CkZquLSYfhwTtSms+e/CVBX5veaQU9
ngMQFfD23pxVLdBkSI3Go9bv+SvmAJCB5Wgq2Ix+fsQqTNQ98eu/mbLWXOYdXqAl
tofLl1pH/7qGb7lLWHXc0WDNt2EXHhxWvIvciDQXE4S64wtVlETS4hubgoChsJlB
9NGoJu2A8tRwm86JSVCIyMypV+eecgSgiWp8lkRptrewJLBge36ZCblQ3t1j7Bcl
S9U8wHXUJS9bA1oSBxBRSZrTIZBqnaxqaAyVZ1xdZ+l/BDcaKp9erUEnyI9MIsfZ
+cr6Q2HtR/iDIsfzPdKjZTqwDUmpltrd8WaG9pmXARZ2Yr+N+AmJw7V9n8eJkaJ3
ntTT9q9c9AThKgPGId9Z7jgw2p0QS6XEdj4SOw9P5hkiDzkIrsa52DLLIX0zK9b2
L+IIkiAjsYl/VwVwqc4bKhhKNqHjihLi89mZUe9DTXSkX003dnHeJhm7Xajg4cs/
GBfoSFZw34jyURJPWl+cnpU3bLmLiFZ3SG4Si3fWsp2SnxRF3qYnO5S0w4IKsqbz
/8XjNvV/4K06lEaZUHnI5hMvMSJpp8tiuIXcwad+Nx44n/IGWsNFBw/ud6WQin45
rj2Nol7h8Xw5YK4ubk7TeIUttgq7mY82nV7MoAPsY5vba6v/l+XLjYeEeO/537NC
zOG2OhgFxgP5WJoUvzh7ZA4yyBF0c0bi261CEWPA4jy6LNrCmZu4tTxaaLFRDTlS
yTht6reXsT42UbDCuRsnrnTmvTgGCgIRMWg////Q3K/6kf9SaOPButkPfxQHMdW1
aHrQaF+HbaTboFB6Py7XXp7Y1wqlo1lDZCC6STbupg6KnM4jEoVMrt68LzhTwz18
QT783DhUuWMUNxwpcAfnxHsgSYkBVkU6d81INvBYUmpZmLtSOaP1LTdUoG/G5bSO
g9n27bV8ghegCV4PQAHSiOIyABN6swSFkQ2ofWV/DZl06zxYdlJ0FhufFgyZ9quF
FuCWqXAejHEyV2yNG6s2uw3c0zwwvSCOX6sxBWWH1wXTub2RKNDM82Tzn3kDSiQY
bcgOm8zIq2X008YSk/QUuhgp5dDDg7vNz7r3xdw7OW+IAWrf/9yQ7Qt6YvZZ/JjA
jx/F2bc7QQ6VH6sjKCj8Rfho503gmA31JgK2o9W2ktjHv7TyXxwHRm+R4rs63IUI
5la4w6J87htZtLBUac22W3U8Tu5vZ5RKy0wk/7YmSBKScxblXe6eMDmFupl9eUAW
8/w1OCwf2gFmaFnFFlcJ56SBSFMNfehKTgYCUbuHDxByWY5YvxEnxsKNCvtF3u31
waC7u2/nTyHCwsuXwKbWd0WtiYRKAyOvHais3BZDK8wZezZXVtZHI4LswCDOMCfo
WrhroCM52AAtXSqd+l8fCyH2LXKM0g2lmB5VNSttsgxl/6Mvddu1VQMs5w1dEs1H
xFiiU05QzmiOujSLmzE1B2W4y1SL7UKkY7iwU3nJ6D4E5GzEItri3xSLt3+z0xRy
iVzcfom8ttuM9ZzTuPrS8k5w//wzWuMv/MvgJkHnOoks2+OSnO2nuC4V3ZMAb1t2
kKSJoB9/VwAy6u5Tk7S1f3gxgG2qdTo8ETLZYOgKEU5aeBMtCoGjppQ4hKORZrYZ
ldUE5n48hCjJy6L7FcMTqavL3QokXGGWfWnIsTJINDFpFlhuDJr1XPXy+uu+8pgz
TyW8cHDFtzUuupN90wLK5KgpvcP8G1Z1mkAxkL/N68RRs+127tSvwv5puopOCY9/
hbu+0GQjoWYNp+edi4KQQvkpKTxQ9zJOVoX2XjnfvPYdqWoo8D2d9sJgcruBe6ys
H1WIhO5kf+CMPSKj8Gpr362KQ0urXHxZe9el98YgZQ7KDl3Nlx1ER1I4wePI1IBt
sS5+aN3O+GLsDu6WW15Ik4Eh/1baaDcWrNdjxvPWTpuYZ8RRrP0P02qh7hbiBlpv
59jqYY3AQW8/yMlX6shQEOfNLYVP29qRgTXG9B+YMuY2PVH2KQ4i3FXmzGPrzkAr
6B7vrCS8BDtzmcCvWLU42HgUwgrG2JHkGsmDkychhijjUHM0ifnMSAFA0p0qLB/0
/bZntu8Kj5C6MKqaimaZ4UXyzvog2rLfpPQKueCCRTbJgH55k+eQZQktzPMFjMyh
VV4leY2unIu4G6rMkSd2FEblLVU2l15cSorBTcjsZ1afpfeBCva+arKcN80166qH
oHmv4soQp0SLEOdX3X8hHzgPXrQuhHxBekPC404nO7pG8i3y6/soA1h/UVPoGER+
e06Da3k9fr7uWpcfx3xKESAWKC2Rd47St+dRSxq51c+PW0F43VfOE/Z+IgeeuFYr
XEJBjhECcNT085ARb+jBcvkjZmrnMd71IyBYz35Ycnlb54ej8AYLt2hAV/to5EbM
nJ10e/xBxmKx38cqIJxY1ORqjKjC9lh6PP+OPBM43WowfopNiGhfY4pdg5+UIUeG
3VJbxbcQd4u4E0sW3bj1Khy0GfyMGV57Tf19bHjk1/mfBi377fINcGECw/mB8eqZ
d5gbS3ooVhWzgayiqPVUi4QwahJMR80QHySwl79B479vapoCmddVNE51mf6BAiAt
stiAFN4Eb/8gsq440qzB2VqgQmiMSy6DgB7nphTHCOeC7/vZWrfgrukw/rFb5Ydr
nxtDJBV+rGnldvD8W/rwiI787PAfe8DyuKBFe74F7bijHGsGdAO5STnEP/6SdQmT
7odud4TchgQrjds7F4nXzRdkDLSRphqkQzIDGYORStsP4SuchKfxaApH9oIgR2h8
7czXp3qxJF3r5OwZ1aKeD8JRMTlqKE57krGAI18qC/g5LfOVxRcTh8WA1+GyaqZ5
m05RGvL2qFEJp0ENo9V0SHWO1632woi7SE+WCqui2p+tcw9f4pz43iF476lS2Y4v
IqQBqbEFP1nAdc4lf+heBoDLh3+pfLFFA/hk1iDH0qMDok0o3oIVHeynjzp4pWRI
ItzprEv8aBtbFIlHHQLsRVNuZeNGNN+u3zUK+qqwLu7MZKooLjAPJZWp/xL19hrI
bPEp2Cf3Cwvt86+1fQDd+9foRjPlHuFDUJNQh+EFtuKbexMOfVli6jSvfLL3JzJj
Ixts8XS/Nu4DVtgsiPC4QaQgji7lD7ZqgAEQfmCbVipCgdn78W/Rnuhtnfh0HcEh
nGq265DBfYEX8ix7YEg7624YkIiRp+auf0nN2V7DUxaA7AIvjZs2eHeQQ9AjeXGT
q+e/7rfvvgVyZ03U9vG9MB6OkmwHppeucRlQrMu1Gw7cWhvK3k0nNenQCSTbP8qE
9WLRI3uknWBQcGLK4MEC0ICNTMf9b3vdHzI73+31RcwGgXJ+f72HhrDhl9dl0MCn
q1DDpYAgPSQiO9psUnbcMbwUvVlc2pqM7f8flu/xtfarKcmKtTPgLl4r6sXRA9V5
ownIRRP26g2vjn7yd9/RbrXkNXY2TYumcK1kSRluGaio5KWWAuG+pO0Bqx6d6jCA
ZW5zZ7FM1L/WTwnGLo6F54pRzgcHLvW/GtREuTER5874MBuxfqufuQqcrDMUYo1Q
CdkuFR6JQw7TOSiRlL0MMLmXlIp2F/Ki/Wjjky1Z2muTkXD67eUyBFpn5lj066Vm
U5TWfqx1Rnq5vj6DnfRFYnP67yQ/Fv7T2HFM3UXcPXdN28O9JPuhujF060yi1Bew
FSjxffn/syVd0hiVDcF00SYHMLlHTdzHK6ZacbKXdPIkZAI+O//0keCpCaraEq/G
KhqRuJEJsWew8yvkVusJNJeL9sYFmYw8yVj3EMD6Kr6R7nXxzqTBzHU2j+Tujiaq
/AaoaNaeVnI9VM5sE8wxkOGtLB+peMIbuDKXPIk323r0TOE0xb5zZKsv41nT/loy
8j+OUifwwXUxzQyBWhyzDvNAdX75/ETIaRYsueyXeO1ZmForQ4bvWVK6j1xThXS1
XHAGzdTUlna6rsuZPm5Am3X2azdv278G4Rs4+fZVziR9klP8MBP5tobQGv9B5u4l
vs1CWWuj99UZ0I/knZY6aUimz8qjCcTd7wTaqpkVPdjS5pl7+Lx1+dD0zu2Q2GxD
ANXZaJ8SrQNuKbiFFix1GBdH7+2SqiXi8QYoaqzqNJXbb0xj0dtkNkRx3w+8odYM
wiRuZkCMF9eH3k5jJ2szvghr2h7pNzRw0jAhq7OMNRqhBf0eG9QS7jPven2o1RII
ieusrM65iNyQLHGNLmvLu3mxwwuVX+PdQmBJ7tpuBwjL3NukJf4jtvrV8JTUR20n
V+yei/k7mPq3FoPtFS52d53dfXDgi0RIJQMjo3y/p8S0BirbPO/CJgL+Bm2WfTMv
YmdJh3o5Lvbq0NSxGGA8GMTbe/8KK2nfqNgPXcRu39bI2GnVricU9gAAIz72rZXd
CYugtagtVKXB5Um4ikuL9kLTqXaFxjba60/JUs+oMhzNgpL70dApHVYijgFeEVyw
r4XazM4+cVCXpFRQ/Jal2nzUiwzJep22gAnJIsEjcGRjasnxaj7F9a2d+4zqJbZZ
XZTG+nfFRWivFX0+AKUzShThGkZf11FG589SGxhKl3L8UFZEAQJg23FAS7EypIR1
95w3wz43fk/26h4dSM35c2i10q0wyLlRtpFwXMJCIfRugjr4Ijej9RG2FJnOFZeu
t0oEoVh5vQEp8KPb8v3EV9sS2ri51gS8MpfOXIspLQ/kEyk+2R3H6gKXBFfpasEN
1Gfvom2iPXU8cWMkMFwdEoYQlgB8QaYOzx6jaNbuyXJFzc2gMNBZKRBMQmxwTEmX
cbEsHA0ABdTmw5FzIeHr7Foh6MfrnSQ2e1w1itE/5keB+3ZerIawBzD4CBVUcOQD
stbz9O4Pzq/scqn9I4FTbj4aqIEdLAQFULBbz3LOUsDwYjvuEmQDhhtjc49fY/44
QYoNvJYidD5JAle7jzjAmn1/AOVz3dD4IRdklSqOodvkBXL8Ih4tYd7X4Feptfm0
ozA7/j+WCnfmkx4pmgrK8JuzAFiXk+1PeoI14zxzi5ykhCB/+rZYdQiztxbvPTTi
PVgqCfPBIaPeZ1zYNmjcOjTRLLAoV/TYF4yqGW9x4qMBpbEGY1cv0ojBZfK1zPyZ
9FoRAWoA8RoZeEbAMGkR+Hk1N1LGeXJXYnP/sq207bSyWe9nZJ3+q2OGEYzqV4Lm
Ziqz+5BCVEeQeSJUdWrs9fYcqWIk3HX3+LmLWWaLYa4Gnw/iJ+Y9YJDOMXUAb662
lt8Kb7xoBBWKnzry706N3/t8ypn4TeGNl6Jlv5HWducYdc/ahEYMTDPzoVIN+CYN
mN0dQeQ3l8CJInDzIiYrzjZEde6LAm85dbKEBAAAr1XADckV26vTHvKbh6HyMVYG
ZRK8CKpx+H54bz5+K1ZUXQHPOXLpkxatnOpWIFVHhCPCldmc5Y4L7DYbAFm/LKTe
u015s/NZviKkSrroq2tbNuIl7Yv5T8MAXTsbBO6ujNg7s08heCYoIpgmmKh7j9JA
FSwKxYFoa8IuLaHdzVsbDehvMmp+plBqfSu73a9hnGbxwlA4eoOqGix6CR0KHjG4
hKKsrCIDWd28+taOvRl4M841EwLdLsOEKEFQ37WfMVo+snfjLCKjfMYelp4m7Meb
rIa7AQUuZrtPR9Vahy7UXGOcCpZ1WxEQtK2WKbI8CEzqNVoNXph+DYop5SmOdYE+
PdLVudXZcCZUtOrizzQyKA0fJJRsPxxjPbRhD99BHxFdn6KAscpzzcHZwmTtUwcf
5hV4MU9iqnPmf+PoIMV3ImR0HGnXHcwIpyJ2PI7XMfU4ibF93i8F31wdpZGmb4T4
X5gDxOiGnuMgwlfGCjx9yk++Dml13+X5EBQx5kwuAJGRRB/F37WqZuc6oyZGffIQ
Ek6Dn8DI+ld0ajB2gxQvJuHjeLD2IczIw7Ahg7NBXgUFb4GXmoaVEVeYVChqhiAF
X7/xtbxiyQ+zVmxPC3KYRU8xWufafaDzDkGWFVgEmXIowL22/CCx0eH/P4c2V6Pv
1NpnnKIO+5rV5xx36euOB+tvLZQ3YK091NmajcF4aH16Y1PTHFfHjbNnRHkG0SwD
gxzypi2kkx6FE7cxSAp3fCcq2AiE8+XtX2VV0/tfBbTEBx9xR+9Oj7rROxhXydn3
UzQJDsE8rsNwIIjLRKDSXSyI657fDxULO+3SyTV2VaSeZ/Ly2oKtycefW7bkNG2o
D/tU4n08/VY029fZRebswMhFJM2k39V8wqDtpwrU22tzsiZNn5izw1OodLMRXaUa
/sH9UKJx3CWXHMzYiWWmC+KqWodTsv/jlkglsiAKy9i98optgKjzqVfaK3h21tk+
/wT/+UFUrdf7dFirazuWWPXTqrLCyNtUIHJVovEQ+fKtNBbzibtyI5sWpsQR+60f
Zv4a59wNqsefBfYYxij/09PSKOHErAb9BdSi9uaeVPLFfS+HFSNuGyhMo4B9/5e5
MXxAbQqoYEh6doS2lAZD5QvlgRWbp/inAfb9S8PGlJSJgF+/GrzrWMGbkSJRqCqo
B/iy8gfQVq6Ol1ZIjugCqst2TxU/ytrH1yS8bBLTHL74SPL81hfdlAx8qGOjOOr0
AKRJf21TMh10vAT2kOSS9PBiznIel4wf29p2Q6+qrBqt1reTOn67qeDNQPoAF9Tp
d3Yx4CfTV/7tx/fmPadblWVO14+ZgYQWwCYpTXofQ36zR9MDwOLaYnW4e9JZpufy
mkc8nDjo5WAJLrTDlmD1jpyEbhWhSDGYcwYh57XmPj9rrl0eFMhN40IoULbR494t
9rvbVKSQUVK5mIpfRaTqeQko6eaeP7ZdiiSM9SmCdcOPv3cxm2OChcWfchvv9vWc
rlwBbAfS+p8Vq4oaQmAXxcK4WhA1UsodG7PzTilh+Gh41SYoOOnaZvleRfzQ6UVh
zJE57s0sENyOOwmk5SQMWqIdGK5X49OugX6ysv/KDamoqPZM/tY9+1zXXX9JhnxP
61NuzVLf6uytpsVZr+TQydFN6rbMNB4Mghn1wQLdBAT739IXFaWngT98FJSHAi0P
JzHxw3WdCGryqegFf+Z9AXXovs6XOobLR23qsbIvGOKQdClm2hRhaksiTfXBwghV
OIFh2GvUDbcufw6bR+0GllvoahsvowDR7GvUeEU25HScwargHBMCR3KtL9z6AWut
OwmpnwUoy+lv7RH1Npf3/jugABo4m0X5G0Tim2nH0e9oXPmruBmOW7+bytgu5/Ld
Bb/XdtPQzaWq6QTMobzsyaRHFNJaRKuZrJV5u4/kpZ6p9s+2gNKvXYOyFZUrEFKK
LBxN8CcNd7+Vay6rg1reievObfCbBElDZQiZYC2VqszpFjYEfKXYEoTPcWr6G+iy
QOBMsfns9kzL54C4UMYQLsi9I8BlmVCfGm7zf4Thk/6pXXCx3FzlKp7U3VctJZAz
vFoHuCN6l6D39aKwE9Ooen0cHR9uL4iNlddSnh8t9Um0psQaOJDljyFbozRjA2Hc
6+Qlu7OTTUG03ruqYRI3PiM6APQ5CE0S0M4z93KsnGlOlzu6QPx72FL3mFz4ZrPt
lr9QxB59WUENr/jlXkVu8zwim7xsAnySjP2SGS+CdC3PfAHw4/trbei4AqB6Iuws
wraDSnHR6s6quCNjX0/1x3JXjFy6EhO6vspG+GGMwlTbfsqNeBGwkkL89ReNO3z6
ryT8ico3VHJh5ceDUpkBeEsfYs6iWtw+hmaH/JNMYEc3HHkaGxoAqX2z0IPNsBRB
4WhnMprUby1KhJp9ZL6TUqdD1Y54FuG+0xYSucdAh0gAtBmZimERT6kjDWW7y9wH
+DCKhTu0LU5LaB2VevFk0SP7g2lgS7gEfJGypSa0bWY5cnYaqxB9AyJ6L4T5q3Z6
oCAzlrW8YSfJid//DoCIEYLkOPjXnbGrjaXSueHKF47y36RgqTrzL3BNai4gsYtK
24XckOvRKcxdpr45GgeRD6DEPJlelyfv5Uc9qox2YPN8vRMg6qhIBZZUh0jrAjFn
5jMM9u62N55qrOWEERt+KOtH1YCC4fg2+5HrL4ynr6hRfhLOm5HCHDwV4Q0hcdFT
M5iqxcvmXFb/BfANo/wYFjVFTxPu6oFqaJszKT4GHfJNFYFdFvQPxz6+ky4i1cDq
Cnw3fiSE13iXHv9DKfPIDmb7q/O5k3zJXI55FrnCex/HnVTILbvQlF7JnE8xXlzr
8i8QLgwPcyp8JljaH/MoZWZxHescB2/F/cVKYvtBI/CASbhSGKV/XYiNq66MSi88
1nTFQg8LgjOnqrbbID7+jHOBNMg4zE96LXl/6QnR3j6GcbHsnKyuUgt+a5Rk3p4O
e2vKX2wODxC1c8xEBBwZWOAbNAGVpR9Q4FxiEZd764F/RBrGLQ/SIJdgzArOYW68
4Zi44NbI3vSeTaMqX1b4KdCvwgWK36kli5edIY6CPbkIp5bojAmjhgN5hlKI+LjF
11TjDzJEUW0fNJDrk5ej5qMmErkxFH4yEL8DIqI5X1lEZYZE2N6D3LekGBE8kxOE
U/pNuxhmy3/5G0SkB+WjyoEcFuXQp7LCgLSuarBF6SX/mW1VscBed5T3Uz62iNQI
03SPd1GekSUSiCJPwne5Pflai3c3HwJU5GaxcfBljqzRMsF6RKd+kLie32oDlxXe
ttA0Ljt2HPOheAchETg4HKWo9nUBu4li1PrIKSYrVdzWLayHnHFlqTGusAIpL8K7
sbfAr2r66ssS3PXOm+cSOOOjugTX81EvS9pggRCbpxWs8RrCPO5+qqbjA0M6MHW8
1Hr2mkjxa659JrjDDAeeJNKAN/qRhm8U6juyjGCh5y+ePPCd7x4E7Nabya7n3oDo
fnuhEouyodSolUxe7j473z+GxHPNDahwAaPl0FMTK+P77htMTenubgMTGslarnDt
aYNgLj6MvM4/LC6JJhW3yJmp6ccBwFqjwx7VmOEJK34NHZVZ0g3+V9WB9Pq2no2V
A68QIzOKa7Rp2REyI5U8V6JSFOtUdvBC17h0tyk9jt1SaWGj8vDs1lA8FBH6jZpA
SY0LaHKkrj+jumFxGuHN3+7uBYlBvyRtxf+CRiP23t4WfzNXTdf0y97wyyLNB5ZK
ydzRp3MMFbn8hQbdV2oQbnB8ryPjTvjeXVk/Eql/wN/Dpd9Mj2j9ka2TwJ+X3+K0
tjCOIsoN6XOG0ntyL9N88vxiwf/+JzBHN42CY7yh1PqPfj5q5PnR6gIZh0mVZ9f7
QjUx1qMYzoWsXWmaRsGeg2W/o4JVz3r7Yu9RE4u0MlD3R1PZLkizkUlKlcKE/hHf
InGols3RBDl53d7YmJH3ypxLK9kJJ+EN0uKO2bRppJQeCtmlxsK1qjRk9HFrZJTB
sjHCsd6zuDbmHLply9hPIB54pipfjHjiFHjF54+aXECq6LcDb3/z0XCnEXNiSqbG
gXK7nBBXjMW1EI+X69TvPW4SvQAERvBI0Q1wNyMYC/qlw8aShPsn22Ob+BvGkN8+
do3k9+CY55LLr+N1+B8QBoeVA0t8tysdEfJakMeWSQbpodCGIbpPc8d1fcOIKXO3
4BIRP7RDpV5qRAx+KXjlbjIJ3BtRAteuRasyvUmu5bEw830ZnKroW0Hwg8HZ84QC
ymardndKdrAw83NeMDF3SpTd5zziuz+3DBZvvObVqEETjLABtHk/SoknNcmUszgd
92tNk+qR7Uz8yFW5puw3G8BwbdN/2LgNXAJRr2Cdsuk8iW+4q/qbfNBg6ebsDoNf
GCjHWyqsGpOIANfDFBpuPZNMxPVYwb+fH3TX1PWvdx/DFYtrfmAnZnzWZGEToq3Z
35TTg3pzazB/aQEgFgdXqyR90j6KeWBFY5iRUfsd+BVhNJkOkBeZ+RsZ7t4OX5UG
Xe8iv6WEZl3OBClAat0s7rHOqK9qVU9snBa9pviFsxn+g99EeyT35t+zyYBfwbIe
4zUhEH0fiWEk4yDBik67KJefNVR0Ueuai1l1yiRL/4TKeIlaBcs96+pyFPy3ns0E
PObl5+baPbcH/GzN8ZpgpYlpsKaB+Iq6KEzyzfWdQGjLloJJUm1czY2MZCsxro7v
mLGES+TwI0OpXymQMw49hODoVB3yTJPASt1h9DJq7dcDD643ZMcDD4jjB825kfKA
SMlVGCJNA5kFDI3ssA/sXnjsKHF/Z7bMuMH+m9S8RuvQKnOzZsX9i61jNDQqpCvw
YNjtu+V4Q2O4j+JPqrsX/y2TsX9As9KlaZTLRq6V6Qtaa3iLL+8sAGsKMg4hXgs+
QjZSBLZ4r9gulsOSY3uWy8/MFqP/dD2fjx0LJe7BH0llFXj3cytWHsKLwGFLn0wQ
E3f2CEhq7CZWmSAvAI5yrxCdhPZfGdq8bvkH8Mjf8NW7uTrh41FHQp9xyvwhY58n
UZAKzxH6Rj4ViDzzJCIc80GvjIkK5Nobu+5eKrw53SfIJ1SM5hPWvzaIfRMHG/NH
uN6W8SUdCC2rfd5XO93QHkkbecJZhhyZSYJc6F1A3BT3IKIfhyFqJ/1XduaGAGA7
39LBCqUMUfws4+itat08IVhykKwD4COeIuS/oFu3NwFeHH9C4voxPQuFLL2Y/S/s
/4oNxaP/Bm1JFfz+9X7jDSXIv4/Tz48ogVYoNjAEidJNv/M9gC9a6IciDA6en7yY
9c4njxvX/zrTTkE1AEGXPceJ5atOaqfuxfkjQIKrzkxAYmDuZQ+eb84wHMGIk5f3
kRi5H22C5YLAEorXI+89t+WkiD2ZwnUgcV1g76PK07hwhqB7C9SE9FUmx9mAuw4n
Dv9lGpiYjpYspwmSzdYXv1itC3c1h64TrPp0t8wxnhGhIMc45tA4ZqmPwMJRFb0A
f5QZalf8tFVgi6dobXQ1FJtld0edtD5jrFr1dZZNZfEBwvEHgG1Z8C4hNCQQilCC
sVKh5BF4IqAtK6syxmOTegv9d56YTp8qcwd7Cmn96mn1vyu9+Lripfs2WyMv8erZ
3skxXZrTvSDvg3/BsrrGMNillMo6Kb2MePt0y1z97yfISyzU4/kE94jD7wt10kjo
uCEvMlDJycfeijehn6rz3iTjlzTd6XH+qIxuM9CLXtyZ44Fpd8QLBGuFOICiTyFV
r8KmYh5zIvUTEfI/EVqoYrvpSMsl4b4GXf2vACr2+oMYVs9FkQ30XwzcmEUEcPlh
XLEyVvQ0EmTtV7rtD//IFk4i8gHFq5SKKh/GNE5dqSDUVJUTZW4NxqHXkVTKAnlk
hwzfX39XgRhDG4/YguuPIkTB9jgnvCQx+zTYny3WUB/2JVU2tyfaio9kePTphfRA
V21frOb8F60LNaqPmiLP0RPsjo2gGVHOuGlYt8kNWTGsfuT3q2RPWCr9XAH3mQN+
TpJxOk7WgD0y2g6sRT2H0biMAtLf9UXFRuO3+xbrEGXDgMA7d38C3aXqonsbV6IU
oCfcgjLERv9nSSBGqAhKkInUsBaGyEGcfZJABRk2hox3PktpOsn+oNXpa5ooZM/+
ZMtX4I8g+j9tOVd6xK1UiO0XD9SXtopBErUuBkb1iNHVIkce8u5Ng5Ki+I/+ISH2
XS8ghfpdeWAIDiqt0drCBiROMkXHq/u/x8JeIMOFvcLVmt9/0A8s2pKhZDsULbJW
vgQTMELntTVrG/C4aPvqanI5bG/u4/fg854Ncj31C3Na/KLYbTAG9JBdSspqJcqE
X2HLeLpZs4ecKW4qaeT0xC5Acs8FMTg89nrJtXu25Y7aV7PUCCjgGCHUJBcwClhs
NRQMnDh7u2HEmrs1arUzlKkoJVyYKTuTV2l9tDKB2F8BkzbgKFpVhoOwGZftp8qc
08rbc2nGyZ49ggQx/Eayt3HdXj+arZwlPfv8zkqfLRdxuuBCongEFPIL6wrXJHBH
/hnt4VFfOoStYcZD7FTVhbn8t1wGGXIdEbvG6qkhdLc1Sanl46IWulOtCrki8Ml7
qkMhWpCnJPlPeGk+6aZq0YJFZWPtNyYYL2Qfu7mHZ7Lh21fBZjb5Wio/BRrqr2Zq
oNwUTeOiZ6p19celU4rqBl7UUYtBGrl+KAue/2cY6ZBt/sVZAw5wKAwTI/dRZ1ZM
U4rEVzZUU1IrRNRZd5JAQarR/Qk3Deq8RZUxvqdEONhfEBsYJuLN6JnzDr1Xv4Si
ZFnAHWvi9yAobSMbJqNsQsfeYFoHl7CkbRfQTpDqPLsj+LwGuKkyo0C4mnhUL3Bj
EQGrqxH0cYvF6EOA6hlBmehYjxjK7AMa7h/EnReyCBET3bVzoN5Kkfn9iZLaWpu1
26Bje0WmzImZFP0rd4BHPO2HuoNd2aasy+MqbLXwAIxDd2XPU7PLaRSrI0eHN+/q
cWoP+LJxLsnBljhuXChtxLHZnSPC+Aaxf6VCVIxqLqAyyBwkTq0Wf3yfDAlkOylk
nvtXbeX/KdO5CLqi8U/bz4pOM16GsHgyq4Wv/hLjiWo91Rb+fQ/yvdMf+iPgYVMc
NNDNzZvyKzRNnsZry/Zdew3JPysGxyDW6RiRQ65hZdlMYXo8Iamo+uHIM5CpBX9L
Hh28Tfwhxb9zr8fBnM+B6UOYbKqOxf2dVYWPqoo6vhToR3s3SW/y2eiNiMyGDxdd
HrGVVDVZqrW4KwOzjQjNvx5IT9CaqxPa04xgXXjqWX+ckEg1nAllGoHgxwRzo7JZ
B282/6Gax+XQpPwJeBFKzlxQC21N8jWP036icHSk5u4Jc8SIWaY1i3zc59bftI0t
yfq+++W//tcYYm3c7HCqdo8alDZMhMc24j9wDchbPUWDShRSCwRTzYxVi+A34TIc
X55QgrIGTz/vqBJuoK7XyExaDIx03xDNPZ9uzF+MdnrKPzaCv2+IXh4L0VJAxykW
LZ4izN3hSN2ewuFdsh6QMGyUvfzNimcfExaXKadGAYRVp9yiSByLwtj/yb+1jjKa
PQAkmLyL58wsdlcZfbVUVtTEpHTm4gy5LMxiec0B2SbUufZvXHvC+0ENThdocDi7
/s8tOrrDzTac6kzXvK9Kv064CvcX/K2RIBREL7lf0JgAlsmSp/QURSHjTPHkurmT
KTp6SnGwImHfqGwirjvkG7vWE2Q68dUSw4CCioTNt3GtFpzeJGFmw5ZnecQqTlAu
1lyLxpJnnVEvwqmWDyIDZrjBhNsKe+5eHxh9VzvK12UVs5oUz2J9dPM/dMAHLIzf
UWLfb0lHRVyxRodTXS1cCND1gncbw4pTwyW5BjY7LEWli5XPMfwVwu2xslcUP7X/
yyTam+YjJwhxCQopJrQlqO+WgwKqVX73eeCqaYnze/a3B2dGx5pXS1Uat6ObG80A
0+li2Fs8uFtn1p3yysek88x5ICE+KqlbTUxezVAAdVt0xotlfEE/UPskH6sXHONB
jzbJ/60GxDu+79q91h3Wk6NsKUkIJxOhVNnjIJX8x4rR/EE69BTOm6H7XRwIdvvz
fK1IAhs6XFy6q7i+2VkHFiwW4W63id4MNOl8Wt93qDToBNXrqJHy5Zm0AB/Mi0bS
EaJfYWE30jKOBRF182rSxbVdw3h2LYzZqV/KVvU1gtjfho35gfHHXb7EDHsvjNW/
ebTBrpsGKF7oCFk68T4QQ0C1zUdCpxF6VA5mXbq+Cj4FhLITKp/6dzCvVJaS3mDZ
9TyjsREsK1QCAe69Pz0/iARLO1wE+ywiFxSh9a0hWXbF5wlHbFU+aqyQDTJiepEo
BEhAc+pv5sjVjlqWBt7mcmIegpahG0feauQ+rnrObADl8Mj1AbxmqGiPWV4pU+M4
p6w8QshLZaC5IRIaWQhanr3T8pa+Q8ainuys3oNBRXlrqTd+v1LJDs0icAs3IrGE
Ckf7KKXiTeM9h4JDRDHfhmeE678+CmTORlfN7Bi1GnEmyIRfXhl7OFac4rhypWYC
zjD0rrwbxfAowvePRCs1XfpY2ECS2EIcTcCVkXZ3zxN+KthkVIWNuc0rNQU7D951
kYsJILo+jnSOv37JcF96rN3HnDucULki0e7SmUH7WZNzkiAV51m8VUHdFYZoKC6c
cclsL4S6XGPEqTi/qSUKbaGAA1MxEslzqQeJ51dt45i2B7UBDkcwSJXI3Wb4MLlF
JBGENzn4q1ThUlJHfT52vvij7HhPYPUXigNfqQWL2Ny6zhbtUdnO3oQ3tA2qgZHI
v0dLvRoYI02RAv7pK7XJsTBPEEG4uvY3swiTHTihl6VIyF80uN3pO4RRHBNLbUJ4
MR0uMJQl911HtcANtlgp9SjUiHS1lDMln/wuTBn6evRDjKj/zRJnrsyOennQ3fta
RilomBQIcVN66t8bu55cS6Elsvp29znanSWbJcqm0PlFYQsf4gbOoBYOjuw5lbXe
lax1WemNVDWaYf9d0WHh46rabwrJhZwnf7m94sxw3ZelfBLjpEyEyMOnHoLaCBxo
AglcOV0mgc0wwdo6NwL4HesBbYGXkJ9P5WnP1nIV7vePUrzUEd2Zo+fpb9Xo5/1C
E/9Wmt3Y99GoegrRdxeHK1+FqG25OafTJARgnsSH5D/itYa3Dq5SOkMjKok1HCqH
6THTZapR/g6Q+E5BjFVap9+tAEMqVdgDgm3FsQ9HHfuMWVPk376JNcayqs7YQnqb
BcqQkiMXH2cngUirBG8whx/VifzDOsUc6ptl02y4X2gdAwoq+B6i63TJo2rivY9t
Gs61CZgrLY4or58njzIwFYWyOSVtwfqbBkiqvp9a2BsFxnu3F/qSYxlaHtJQNa09
CmAhsv2Hwf1Qi9w760Y92ZBf2GzHCVrqWXv54XbLbGUwKVxt1qm1NlQaugvvSH9F
/NSBZz0Jfv/TJYZq68Wsyu+CP7u0i1DR8KJKTStiEaJ6nHBIa+76GjK5/k+EWvk6
KgFREarOEYDtbU/Vsvy7zuAAt8IC0B907dK05+lAFtMFomYnWryDz457uU6uHVCx
ZyM+S8aDPKzQhkc5L9aX3UGV4rLXP03RtStE+9RKRFgEmzsWS/0Aww/XZoRbbDEt
fw6eixdbBe855bLPQcCRzH35alUgKngGcQV3ZlYro2QxlxV8bw/T26mcna95DNqQ
T7fksNLAhmBYRYD0q/ZijsY8v3X1RRPerKP0fmGm7penIirO1xZ6eti68J8qey+i
Y4mC/MYTSe0WYoisMT5e81syUFbnby5wMXy88lDhvTjQMzfqFd1LnaB+RhRmrXtX
qMW0gA1HsDSJ/WyD9puuWI28DLcHeHS3tkMB5L85LYvgNI/HWEStNa7StQ7kTedI
CDDpsXQnlN4VGX+oGdJqIB3yGD24ObmMmpPMYpB/QZCwUiwP0XiEvcgnAZWERKv0
+6VvYAOazX+xUPB1cZCUx+hMmsSCsGzEPLKyhlKuLeWD6W78Z0iN+oJKEIz4Qdxr
2qzdyFQ0fbMKuvTpMgGfNhR0cba0RpaAIlkeEQdlCk+5TA4aKa+YuBhtMjJnkr7l
RX/2miLol//3tPYi/n8z2Bd00CxRRs5qYxr08946gW+dX22MUflx2+yyEcCJoOEY
GImN6pk0e2E3bE2nZwawz0Q+vyWUUNzK/9V6z6xu+1XYImqkvJsNKNmmhvjJ8CL4
iPG2eKfkNa14EX2i8Mcz6o3jML/2N2wzgQ+WMa2ce5vzxOQQ/DRfXTqb+QhMMNGJ
bhe58elBtKE4AVYhR60bZc6kSchpRhU9qvJhD1Br2INZT/t5KGYmg0I8WpHHhziK
p04B7Y/470wyGe7vmH0/jA3KxtoPaTHgoKTY7YUIIVRSE6KSj5Q1B8Md0/RrlVR6
yV/p0Okivli3tBu/aSqD4ZUFkFdd0DL1dv1KlpPQuZhJxl7G7Spe4JyU1HtVv6Ey
F48zVGo+W91Q5JTcCyQaVs5Tt4Akt2AFEFRnXJwAS62lLUTiJ6jUeIOEMiE0txJh
9O/tS/oVzd5dltpFMyQzqEypu0mT6poxfcdqvLw6YjS0OOgBJ8OQ3C5TQeEDwU3k
FoLpv/K3vvZoGTnYekg1vDE9JPmCfJrkgF/PhK3jlrbONLk16dt4Qg0RN/IN0tMh
pcIemTEykmZLXYxAJ6UEXQrjv60/dzU1q6dRrhv2GLJh0LBGZumzTjibN0cZdddB
myOY0Ipck7OMN907PiqEG6Q1zDuYKKW5sh4dCWYysVFLMH9vG5YgsOXkKbsLjS51
NSs1A4AiKLrOW6POMX0YAt4vbH184Q6LPnC3T5oyNwJNDR2pbmeqCO8obnubhCi4
VwzCaT1Ditdp26dNeOJLnAxHD27tKjCpZG06DTm/r6M2hCVNmjbHPyva7t1drJ1J
Jb5LRN46hvcDhAO/zn0Dkg+vXkIYOwE311neJkL5A3XaOZ1LeaLCUeEbWvRah0l4
7tTo9icMkw8ZddDcl/bLlsD3sP051n8CnMiGt9Q/tGkblJHWEC/Hy7OJ+gP5exY4
0YmtLjpmc9pTS5qpWdu5pLN/PHaPyIbVhy4a5oIjM3v1BdFb9i52OsiiYAn3iq+D
uuZuAEy09QcgsFfMJCX7TiJL5jkJBmkYNX+eHLcqYgb33SVr/1Ipj68OojN+lGAJ
UpC9kyvQmGBwDnc5oSvYpFV2f+M82aL4sg6T9P/w3mWBz1xjQaYzrK7NuXpi1vd8
tPhd9A7EV9pK/ZyaKgaJq6eNkyH99BpwFruglst3HXlo6Oytwpio6W+enPyh9YJO
rWjzHd1fQINZ5QHv8p+2u+krIPcUeZXuhkGy3KpGEIM94MvizKOSSbY9qz+mmOJ0
FC++WRVCvR/IX8rp36Fafgth49Y8GwPTDPtOwB9/y9IHyDC/YRSzcsVQGVbOYgWV
G9THN+36HlofoBxAtHCncMnFJvMVmazS21vDZSxo1dUWsUxwLvYtblsCi/j9fCix
KKON8vLXDxEEES0iMDQdVYlTCAkLBvZqlwQ/ujIaiiIDBwkVwAxHU5p+RBnuuH+q
2f/3Phgi1B383BcUtl0dZA3cBsWPoaE8RKVSgcprSsdS7s/ucO6GBAOesJ5fbOmY
NIjFmJn6RP5fkDqWQgcHza8mh5tFcibbG77awEGeJPCBiLuecuQ1W+FQk5uHZDTy
Cs0ixPqW97RUw3r1zdhlArtnjSxkxfd+jCSQtGMlj80VXFjSN1AHcRxdCyYd4Pl0
lNq4KyO3+v8kB9H3cXmaEZtfbThUQzb4fPx83vVsw0P1OTOyehj7K0YNm2IBh56C
6Vbkp4k7Br9eeOFt1ltO/2qQHlH2e/z7jXrsH7CXks77j8owRN+a6A1palo1RqQS
USIoayQ7v3riUax2nfO0VSt84vPBOWCYux/DSnT/Wth+ZukuB/YyLAp6ouIsePW7
pwJpFJ431Atxr3a47/sjlZamGleqFyxmrEnSAsi67RhZTkyv4cR52X3BT1noO9IQ
iCuSMUmm1VBd//aX6M9YZHEeK0/WpPQTXtFLyBE2lMba1W+y8MjHZf4UCaPu6GBH
T3AuOY3bCC683Uc7kIod/OGfYsJcmibrsc9DimnGRT/2cVlln1/MjpS2xGY5Twgp
4fQ4AW3ybOg2A9uelZgqGCx5a+qnMMAlTrXl9YRlbApdOcsTmWxXeK2TOf+yT3XN
7Z4srnieb5UBQjKcN3JG6AYw74IbYqwysrxfE0AGTQ5dJmuuQaoZXgNS0A6B188e
J6WhIDwLgqNd3iKP6rX95QEhFaXAEM+GvQFLEuOp2FFVA19hVx4fUywhMnBz+HNi
ngTYJzgKq5Lm6CgHJY+ugWpMdfl6ZXOoOse1VyM2VGavrK602VzEPG2elOsHWsTl
zRTuIMsz3TscIv6dJXIX546u+6ja0wTmJvA49SvVougvMg+XveOzRKWDaCQAWBIR
8IyDT+D4zrao+c24FMA80uKfOLnQgB6F4s7hQj8TWxVNafRXVExbfySm50YObYrO
zGqgffJpnmldMlOEL/vzxZsEFBxjs03bBeWMnr26z68siWnOx4Ci3ycBK6T4xb9C
FT8fyoCIyvw0kTREAQCZa1K99swYkDxCrRz3MNRuf4vpRlYVknQocP3nxVBQDOMR
aPhNTMB9nWUMG4/NqcE2Zn+1yIY+dJLsDC0sSkHYXRbX2Or2n6K2oAjSSdfiW3Jf
Cwm6bxyp80boyIt62rsOtpCA4TXohe8s9ijHlegHuLqvKq8auitSsN8KlvSuOgJh
Nk68qn9uLqwXEdhxxkJjAntAMYkIKkDMPQSZ2Ohn3k4WeY/1U0ZvcKDxzLo2P3V2
Ppk8+MIq6rqaxDKRPfws8HAJHqOtJ3ozs3SvyZyYxlndjSglgYfCrgpBX+3vjeE0
9nkmifb+hgs63BltMpRSDRqjJPdaaL5g3rQ2Ou3e1W2+vbP9uONFAAkbhYm8YFbq
cygLUgrV7v+IwP1Q7f3MdDt4bMikmoEz8hH2tXV8hpdW9mq1mtG3WRGjjK6hpZr7
NfCawmyBOZej0oKWpokccz3z+D1pJHZFsnqgcAnZgnw1cmGhjShiTn2hlo/5SWON
bOsQHL/xTX7II7TeoGNMEaHEjIvB/L7gXpDsTEoQwHosVSz7Lc4gFrPZouMlTkfG
Oh6oaxgfC2VBx7McIzi0FCjX6oMaw+Hg5mAU558fG5xghXHBClmbr19zvaZuDFs3
EM7Q3sXDz5Lv08h67COuiMq7nPgopaaSeTfNKX2AT0MSI7PW+uiE0i2KwwhQWYBg
WOOEEb/rqPMdbPp3u4aY3JDCCSAakjQzuK6wtDFw3muZllMmzQAotCXYZNN14LmI
QTVTXSCKjcNRKDS/5kcwdXgKlq65lcNjq0mx2dt8ZJk1Jg9aT5M2ut/MWxfJ84Gx
vz2Cz4+BNJkAmQD51wNGZr0ZJhA6xZALTFulWoonM8Yic7V+a/ceudsHB+smMt1M
Ak1rUf0tcol9gWBg15ursWyPurxVfCl/RY72CTFoABelpKeG8iCswh48y0KffL4T
Y4kkuf4xWs2FFniWY5d+jarPtDu0QRb0+l+AWrA4u3huwFUV+RpoyE8vPHztaxtJ
jqicWeYRCtaUHnMIOD6YR/xMhwBcyYKGY5LDxTxujQ59vQae/5BkjHFY1oXwmjHu
CUaiOdivjfL+CHMZJSFpkh44fYkq9UXSOjmNNKenQHBjxP/xlExtyRE/lyO45XGD
DKE5u1v3/O9yVu0LkEl/x3nobj5HXwt4zy3N7lz8bnxbe7IuIupbbj0r9lAAQ6qW
JyJm8ZRkwhzGtLk+1+Vh+RVbcZpUq43/6OmvC/l+sv99Dcvl+TPzV0cf8gZGJ/Wg
QimjVB8Ax9Xk2pft0XPXJiV30T4c9GjT5gCw12SEPyve819xKdmVws4etH0vMbcH
f/UtBfvpj7NTsBF6SG0ZFCcmgkXPPtkFQZKfuj4cNX3ep5EC5NPTshFHAFXWUdAq
bFpRp3Tm1dbyaTBV499XfFtnF6w4jtQprMUmXR9Kx/zZJ6BcBvL4dZ0pp6Hb6bth
BFct4kDLfKDZBV+2rEbEnhXu+4XPW0N53oqx4OeGGUZUwuDJNVKUoCSY9tPH7b/w
ujaib0sruT8MfMKw1ooW5HF52TrxpA5a67yIgMtkDYR7GDgMEB+jL4PR3x+58qNQ
HzG5PSaVE3677v9YzfLNIP3uEfAnqO5U0ZZzyeOT1rf/na80DU4Y8POo0/dreavG
KyCIbZW+L9H3a4diXNAYVZuVIaeqzz64GcXmfxXOXLFq4gTaveNzXHj2pIWuG7kR
JfM9ivPl1fjeHQGJmK7vTcGlxnVi/hUxMQtD6aqYac4GIyqK7ZfCa2MR3zgUbtBi
jnQPbyXMHw/zj4a3NCwTnwt6wEOk6bYNrI3oNTaa+TrUNlEVjiNSTSN/xHJn46f0
+6AE9cHHqskEtst4+GsnckTmpuXMMw2iECQ0YpsrqtY2osvnoHBmw4Xjvn4VM/H3
HSgl5m6VjaUYerjOwMbTBezp7dLRCerd2ERrPc9gFBEMpFgU77HmlgFtU4mClyAL
blMmQ7KIZ9A8VsZVvqkhgUzsXRzANRSOWoNUdODVPp0053bNDxIzb1Q5X5rw0WGE
jbzlq12mj/QQuiEaPsvBW/NmFzsBEMG0hP1xdsQJfH0x6tSTGYuzv0obm6/IpyZW
YVXZN1hPto490/5d5gD6gcjWELUii2UjhRdPAKwbqmw9BfmSRpwn1pdgC2l3iU7d
fP2fNBjktUkzLmFFgMkp64KSHRVeK4R62WOI6x+pdAGXjPtWRF0xfwvlvS0j6G/t
3vSLO85j5KvtqQK0MMvK+1Qez1/YZzDqNYy+xB4WfWLUN6oHGTNBpuuo6j25vkjw
TtKMr6+eH+Qd9KirlQI5ljwOYlMFYzurBcLtr4hcbOzSubECiOuFh3Hk4FOQktp7
+aTKPACY34j8btW6XYNG1Zne417zpdwxvBxJu9Ugba9vnPLLaxVuA5eNjkDuAhNU
FR5CS+qfDBkjVzBBxRj1UPW4tK3c9mwH2cpAQa1Lrc6iMzFMt6ewmKlKIDCyPrFf
f7at5e5P3q6pFfwQGeTacmQxQlaC9KZLZPv8ZITArGZOipy11ne5Cki4Im8Iy/bJ
czGYSYiCnJldr00fnbuEQvuVJyO9VE4rx4d794AnA6KjkrYk6M8QRJOY2XNbeNSZ
uCCD2iUwhGHGsk/uzp6Y3UG2EabNKYOAfeFzqUpBwx6vPpDlfy7n5SDhVcXL8k+o
f9k9ymKOSWZii+zhIYvPF9wuFVSSov3ucVRbHo2MqOrFo9jRx80OT+I5rh8YA2N6
jGQSdfXjDhlvNFh+mGXbJIBuDQmJu8VTaMjR0aFAyTiAo8OKyeR+SOK2hUs2+mSo
OaskAOoqi621lquzDOHjehfkOZIeudeIbYSeWSZTzVCYdp1zVNy8MM6y1L15OZEQ
FwmcCsq9nt1jUy6R9zGKcnOftN+s8H78j5aKjEfxPw+2i0X0CC3UmV/KcbFVmOHN
bzni9PszfqwEPVALf34Esh/qJ1Hpp50nPK7ZEmOxM6DQl4Nffjdsm3WwK5XVyvk6
7aNrYoDW+kYmDU41Jkc/tgEYeITNVVSvlBwBHFa00NChcMXWu4MIjduKcEQQr+wL
qkw/irBAv/RdZBQstolwNkDIE63SskUqMo06TPAb0jk7YrHq86wDv1KYnnRI/7Md
jFMCes3Rrv+xiNuG7ora+W3FogvpmXhMrA0+jdURGumyM/v3rYu6Kuhds7I+qCm8
IQaeP3E5Ktxjxyk6DdKNQUNbLzwuPQ1UjZmU0fnW8Lo1mGCiKke4v8SqosJbT3gn
huKq5fFrApMzEDg8IoELOqXqnA/U++8NbyfOUGUPhGKY1/8DML4BoNMR54COJy+g
aXjurkRhQDI5UKT5JFt9nslnoOSWcgQd9XuoRCjM8yYib/NPwjKL0AXwMd+RjeSf
FWPrrPzQUq1Y8Fw30AnA3DPHOkg2mOBmRSlmtPpy5mTQJuCCtYcGGY6Bitcds/D4
hJfDvcwU/xrPdqyqJY15aXJytC/NJO7WQ1nF9YvwraTThBd+4H8c985caQBa2dGR
Q00sGkZbFGLQo02mqW4ybcRuxbhYIfEBaGYZ0i7/o5tV7PNnovBnVVDP2BueqsJx
s/MbOie7/9V2opBbkaMve7qTRTxH0aQvpqlzcDHHuqdk1/PQ7C+qFz2t/Wq115Ur
/fAmay83Val5fniRsd2dOx3XLrB4nAjDbZG4+Dr2Zo8atdHG3ubCrf/IePRidXPQ
7cin6BeKACLnfyNuIEzx98/XPnO9KSjImwMM9MjXxf31QfR2amBvgPR8Lj2yKAQx
CcuHQew8A9CPSh5RjRBU+14LpYvSzlZGcPxtpcO21ReO380uJhoKoJTcdsFaSjUW
wu7gPTKDruq3CuiCYGpwwxlmI+3NowTae+DXCs7F55HQU8qMenucBB6bxzMD5+UD
dbtFArTK1C3cuXmAeGN/Ng5DSSglKCf0i9Jm3g4v0whoCHQ6ZyWyb2x1NzQlw6RW
FjNSzurO26kkUlSy4+y9HMEyooWnx5cVTUGtljUnNofdn0kODSm9AoUMDNNFpw+g
zGTleMp6wQsdtivtec5H/W3bnW3O847Wp1DdncWZcdDxcNDBlLgA5Kc3i6v++ZgK
BJQsv+Z01LYWbdukQ6d+G56hG4iy+bBpwGkXQZftaU2AZlMIRVX75qzaI+FNiVvS
sA938f1XwLt+S0BIOcuGZWCNTCw5E/Qkw0mLbQZVmHTCcubgGosL9L+o9PaKu+7O
dthxrG42LFgrDMG5LixWlgZlrxeZ9NAVJB6TSz8Mawas+THNIyGMFnBpawhVGHz/
b83aBLpvr4Ltl+SgkhRfoiD1pu2RsRmyBKSyfeml4igqr0KJvMvrvuizFpA9JvsR
3XVw6IdyS0mF5t2ncNTZPvc/pZ8ECKCN7Qlp7+i3DldL8WRgdiTvXgsVQN3D7Pm/
16i/Qfis6mNIy22E3dySVOZApb17x+GCaHJ7/sVV7oWUw9ATyjKPjC/5Hgh5/y4M
g+YTWjV2sUkCAZ8ioyBnVMajvJ2Uos0HXHZ0ZV94HJN/boA5dmgSXY4CIXybph21
9DapHxiK1AL5OEu9cUTpoQ+i4gcUKzVKJ7ke658Osz7imaR4pdDqQhTq+cgiJY9E
NPuzfCb+Yk/3m8F4d1jaF+DMwm1TEdleJ8ca12nNIjarV4kBPxpQxK4eGze8Cj12
QOXkE8MpCfHgvleejtnngc8kihknr5IQFzJz29eWdS5hEnPxhw4qV9Hsf0Kp3t2a
R9iFwoEWn+qtzi76zE0Vy+ZDAvb6LFSEbhLhOIEGtlxAW5L/5aJs7sJb4sv9rKNZ
CA/M+fXOuhpAG+f5kOi4wSNFrP7YuUM1wKFnBaa6hOveBxyIGZ8Y4tSr+TALWDLt
+CRb3n3W1rMXr7foV8SagtDTN8cFcQC/5Hz6+i78+GTZNkmBgnuQXNu5mlVqUWmq
CPi8fgSZKVi95EM7eh8n3XG2bbgV0y9DNbMhmNIl0gag2DP4blMKa0rnp1npilu7
Zb44cGnZkzrlOfZMfYZgddkYtrAnVkAcd8/W42o2bYdSsPX4j1w0O8+H7h+53Qwx
ZlEb/1Wz6A0mYN5nFhVZTI1i8LUNZPl8/GT7N/nsoxdpivUMPTwkEQy67uAhExK5
nCcTDcW3Iid50UvGvxa4cmUGuB4xCiya/7Rq9sK9qo6tD1o/LjndKSBSmqgVwm5S
WKCJJYlDOyR6zbjkgXwQpL+XEYN5sy0CnOFJMTwZPiLw3V0SKZ0Td4PvzU2e9fra
wh94WmcykLx1VkFY+Ad1chgXSC9nMgelqwa04rO33yg64CmV0xBlZLcjrJQ4iR5m
hd2UPwFA1kIDSuxDiBofmUSHjSNsDX/PbTPMH6RuiM03M73GvaqM0IPm6AsvEOh9
ZTEEWcG9XPAffKVO+dqRRrmm5b7FGwd7RA3mDUKGKD6kQ3/OR5r/QeELJhaY9j+z
yBzLp04eD8dqugtyp7+hhnvG3WOoa4fuh3Ozu59igPVpY9MptVJoncfj26di/4Q4
taU+HsKaaTJgqWwQcvIWYyrA2vbKpBCBQHVC+As6Gtq8PdAqzOq23ftZxZFiokq9
XsZ4k9bTCcuMqUSESnXof87/dv15eVOa2qTS48t3L0aQS1bpgj4UcJhj3hYuDqVI
G+bp7eJahhy246Txbk0K99hfEmXoTVOW7tP3Pn4Zk8G0E9kK98/GcLuVnozzaSHB
YPV4d7Pr/+oTwzPSbFcFscIM8cG6xOV5LXQSww7jVgTZuA96DAh65p7WceYrX5JG
2Y15JH5iRc63kQy0sOt+l+DAzBeicNCkamAHOMuQ1r5RyK/OabzqGZvyo/HguAkU
TU0AhNH23ztAvGLYuDR79wiX4yljY7BoPXNFjjMA9isWcnyE/+AVpDkd9mCIxzzC
SkgJNSuuxgAGXSybDgKYDpg8KmDPNlOrXCHu0Eu78zkAaOHGUI31iJrtUUh56o2p
+n9qvzGBr0HY39pspdZOtZqC76V9Le4PqqC32DWbzzVZ3ycoQ7wElOvppV5w8kEt
zsTJLc2q3YWrn9YQExmq9OfsbAbbdNF7DuvLrntY0jD0K4f7fwDGvfXhhAAZnZJc
h/IlmXEgS5Z2arrOaJYevNikRwkbuzDW/zZm2HRtpoAlEGN5XGSSKXb6b1FY/Aye
9XTwrClBWrikjPilS90kVT/nBxZYRwrcfxAMh7yLBx5xsL2TRYSLanx7UQZ2r9fh
qeiZv6SHZTayJP6YHO0TLgzeJUEzhvt9f2mw8xn5H07KkNGoEsEUtJxKyk7fJR5R
vs7+dpI1uXcB0wSSciDKCkbTxXErjJ+j7CoM4tCA5aO4Xxbd1aQZgPGb2g1EqOfW
1pBBxuyYHmW1gdARCThIokChwzLYR/0Y0eVjINWqPZxvmDmN1Kzv8BAC9rTscgeQ
r/yvDW1FHAaJoBN0KXB1XBgNo3XhwagEINYkeAbdGJKHTLRUhccYtiGoFfsXKOV0
nf+Hjw7w7dXAh+YUmXqAkP8RAFkQdIRYqdhZF/RpNz5FrO8gk7U5P+Vz1RDWhmnO
L0yUdA4KMX9748tFSCNwZTOH8sXbDvCoKP515njHL8wi/jgPiojbENPTnK4Dnnzd
W6gSk0e3CAJ2R6GXH3Fuae6LNcp7Z/kg0msvS2aKXW+x8mdi0+LeA+2Epb3U+K22
gMZJVg2Gv2rdig/1SzTBXcv5tIOKFc+wmp7OYW86U1XZwlGaHP11aSAff2G1URhC
NYINqBIWEElw6tDEWNOhxsCEaX+IzIz6DR2aLfwTHpZ2RjR542iaA5sHnM+YYuz/
XX08yNj0K8hT6RPJDiRVpoajkT3kbAMUCNAry08akX1bD3g5zB9YWZscDpKpVbLV
HWaF5I9gT1wY4cK6zg3zRMpNyzPqj7W9JW3w9g9KlWY3GEOUWjrn69JcenldDE8p
QCSPIYP73guNUsLt5zljNvsJA93Qwp11uv70eQhbB1766p7bkD7HHuNRcB5od7Ah
lLMnSn2Q+m0Ss49FUlf1Vk+3igrC6pM36aFARZJ6rx7AZlw6G16/AyVauJn/S3xp
8CwA1TPn92OYYLeVK2eDdUfO6hyXdtfssxJntV5GKR4tUN/Mzd19MS86xKFZgpwp
Pou1KXzsfwnySdFj9q5xpKnwZ5s2CWe/0h/CFaweTIoHyt6j1sNvrtNYrDi4fmHx
kzS2k1ErQCWbaqbUyXCc6i1y9RTsLcSTAZkic2sZDXce7aDVNP1PKLJJkFOXEjXz
J9Vc5P/p+DuFNeDEs7Zs5wOeU+ScEMIuliV8mGVAO9iFI9d5u64TqyTQQSdK3g+0
vxn5Xinn/0/djSW3rVyTskmSc/cu/Vj+kSZY2gDpqVNLP0Fv15VAT7/VGdha8eDs
EKKchEDs0USbTtUrQUJnI1lwPam3swdHASG2skjawMx4caj3jqNF9hirfIn+FOx/
iWfjzThf7e9vTR6gvjFH+2XF6kDafE6fBd3+pb6b73uJMamY2p2gNohNYgEljVMW
x/D7Pb2Da+OVsvuwktuK4xudyCZVazUkn1FjojUY9o9tXbIgchlYOaZP3CP5AeMu
Iezmfe012b+o/t5ejMH2xnsi+KfjpYNyOsifkPHYcYQ83Du7hZvzd1R/XESfnySj
t2KiaJy8dUmJ6+YQq1tJYVMU5N2ecbRyanU0zVoiGW/CQZ+4U4dLw3g5dKsfSCnH
Gbzuo0VG1pKyJsgaOMQ6zRWUDSDGeejifzLAb2TmTtZiQGxoQONgkS/wVi2kSuh/
BKHvJ7Nt198+1TjX5UfdC8VDeVVOKQEsDFbE5/WL2uC+f6TXutkAzSL7ZIoLy6zr
5QsO+otQjTF3H+ISxGfkD3KQ39y6FGL7raBwIQF7kcUqKlkDFUtRNunGebC7Xro+
jrMh7HSMVSb4ViecSVocoEPG/LIfwO/osdSjhSX8kxVJ2F4lHli+PrL+acE9VCAP
mzgNhib0lmBoR2hlE7yFV84bljOnRheNpWbL6/borh8peSfK+amK5++lltdrTs6+
sROcPt+i72nbnyhk+T+1baZexhlslh5LzZgTVbT22zQSZ4bkciPEKnNRexqZ/sV1
GNxSj4rqhvzSyYy+BmQ3x2AIcuHwkx3c8b0cbn9yrR0O8XtQ2aoU/6gulxeNOMam
mj5IyepD/k8M/sgF76dxhcRSz/FO++p1fRC4eDA+EnYsNl2SMvNmcdMSRO3Hu+PN
fIsqkPh5JA9vygB+0X/PtOko+vnMMSwlOvjTrUlhEFvvTtOZHzXTzPa5QVGWAvX+
eFZPeiKTv2JUD3K2p99rE2QlYSG9rsj8gYDwEoCMAIXO13NWp9aD4Za+d117dQcQ
h5x/pYucrH1le0D387aIbus1oaPkKq0VpQ9obclYC0YuezGy37pbfA41hRDGDdY4
XzU8F2YLXNdAiWfF0nf8fdWVtzcgrdDGpb9wHvtw6PpRekI3P0ASoh7Z6Pxjug9h
pf3hGt7RTIdkzze2NgMFTbIEt3nJplGely0el6+ubi0JHOZuaet7Ur7cSAvvbxZ2
54PLdn73xJDl7UWHHqvF++AW3SzrwD+a9jdP7U6TrE23REWq3/X+opNFeKpDHv2F
4C1ePKmCittoXVwytGTXpO+4E/dUt/j+FO4v0G7V4T67jTSzksGLYNvrEdoEypFp
XNQhLiMvF5JSXroE257Dr2JE0oT9i/nzZ8cdASmfzwDyjiXPCysTdIsCltDIYJv+
D1HCY5rvWdoDhXmkiB2KP6sO4N92qN2r3rgxpXzxwtUZKZkZ2c7VwwmV5Sb4gEVK
K7DNP1uSrmOzSRgDki1iPuo99O4sxi9Aqy7oDwJafA1IOgC2B4y0D0co7WgdutaJ
ba9LWNmoNzp+LssR+4Kof0Qe/ia5RXd5rXzLDs3vNmDm40KXHuZmVBbnU6DAlEL3
XRSPniB39jV6W/rAqOqCWrmcGxHY9GMV6IeYiKONtZNOABl4YC8qCeqZKf772ZKt
P3MaWUwXuNvqqJBqxlmzaNepZhs5wBOa/zXROHbV0FqGky2s90QbvlLsv32KOO8B
cDjAjz1KI72x6RKrgduQuMvEVfVukRayzbKt13IQ7VnJ845ErCFO/+AvUOkbsGI8
Wgi30iwJBCAGwz0Dc1ehR3JhD1NkiU/ROJJGEoOgO5w6WqhXRGpHsxc92Qxra1AW
qlL0zS/StLKaWXBEReXDAhuFRYCWG48JXOAVcArFtjmEblsxuA9iaUyvy4uqrQsx
tvznkbmtCZ3ZBx9qcbv0Q6/w8ZmENYGLCp7SER3VCFCwL05VwuIodYiy6hMS7DRf
Xjx5O/O6nY3L1Uf48SwOtq7u89L6jmCwarqHT5lZPQtfOhHtAwENc8h6X1g5PgUY
cvS6fxLiL5ttXwVtvmKKKxjyqiOnixio7MmYViBFZlrOF1bvOaYgZ925A9qwBCT0
35/28pUTaX+hdHkE5L725rv6b1e6uq2SaHXQDk4dXP53zZZSLFvIsYJvDgqVzFnL
0wCyZwdc3vwr6aU4blSlexV9KuV9/UuTas1p+DxWL8QhWn7Jky+f3Qb7VHuXIO5W
r6v1sXzBUpkPeZ6vu7bCOfgVslKQOiD5pWU3WD4VWk3PJKlVVBfaEv37jqqF5/DC
60aFtKw/5RpbiPF0QEfBNmWxmN1FnyiO7nERHFnopa1I0URo/ax4SJuC92j5bidP
WrvJLMLaMkU7Dck3DuyOP0FxH4RqapJ/vWvz/R04h6hpqhm676k6bVJCTtL6yQpS
MoioqlDQ10tI4B+MZE9WmQCV9HRmAxprJKhTjJVtgeSyGzXpPG+rV8ObAnSXM023
PXlnUdkE0eWN7a/OaruNgE3wQso1uHIP6cKtLmU/su06eZW+FDcNC0lSV80/XvkZ
pJ+mDrlkZ7+Do8xdaE/yGtLiT7XJC6aJ619W1uI3BwjUHC8iRu8pZuvQc3/b1NZ0
rmfI18snGHX7IbdVhMg1Sknzcm1YJc1SmZkTje0CdnjJH52VDDnTGxqtaijVyqCW
SdYoshMX/ME3dH5eIs9g2MRYl5rSRW/OI6BOXJY8uBJv/Sl19CnEhLgEFQ1gViaf
5l7D4ft2ASFPfiXfkJnv+zWOOdiynlfJGoy3TOXeRO2S0bZQHklnk7I4RbLbQaDf
BglUMqyv9lBYYCiDPgCQ12rI9BKTmomdz5qtrsCMVz+p2t4dIfmeIativNbjcHAt
QGhacJlJHBEQGF8gw51y4KDMUt/rHGWOY5B3+JFOJ343NqoZVsKSaQqEePPxQsZl
FREeJT2GuNyhn8+ueCOPaBSubNiNDPlJk8DqqmR/3Mt3XughHOsmxdrvvfjISeDc
N7Y1hMr/+aq1xrojye1JJnAMjSpy8vKLWCaL7kbw7Qtg72AZGFf0w5N1sEIHsoqS
cO1q5Fowzczu2luMdGTa+YKLluxetiWRLCq9u0FQNYBCiJX1iZRX5wXBpkVGK10E
n0CtwIjaBM3IyYylU13DNSiCxuglX9Aj/STvntNCmolAwrQPIi/srhvLqZWgHGP/
Q4jvSzu2R0534BihLPEznPEbA2lUrLC6rpvGdD9PQUvTO7ekvZhbV3kW5AdJ75j8
SK+zYw1JvlGjjXzd+G4ZzVW7rE4oVyleuz6RHN5ZJlgurEb/2Ejp29mUjUvVSdkJ
pwU2XQIetU6EMPKMu5tYeWkKzXjtARFVHsV42daTcKDJQoBgk9KFqCdXRA1WtyjY
wqYmQF/7YgDsWOCgBffSrRQS2pukiHY4M5+D7FB2Qq0d3Ba1XKks6ObBeQNBjrgp
FAE0N5Y/EyEULToJtpblpr68z+lhs4v6+W0VDhN+GluPkWCz6gMzoF2p1Sq6hbTm
dbtlJfozY3CbtEp3WmTpNYrHLrbS9162H82joG3PLCtqv2pMa/Ew1VyJC1hSQhA7
cxNukvnwHt2TcxDjc3gBcBLS0laj6bekJgB7RUTMnV8YI61vU+3a++szgNFINtjr
RBa229p/Gm9jQM3Z69vUV3Q5XE69mL7m7oLhFCWzSMuSSTg7XXS/OT/+QdrtmEXy
zdlxJ8fMT5N/Z7ius18VpMSGQRz//jLidb/sbXnF3Wufg8iyniztDgFc1M4B6FWL
88nqsUKfhn0ys5jZjUJ8EZn3z47nJd6S2TFuKL5ml69HZ533apTlNqfsVhJmAaH5
18UyTktacAxgo8IcAHICZ9PyRSi73qE5qdpXk8hQtKI7YEiipIeUM2dJP4lPpSdC
2xOgId928UzaDEXLArziM+AVCyobtGbDbIoH3+LOC3RyITiKnX/QmhbW7vIHZU+P
cwNM7HJu5xpyhsSQ3Qprg3fLZnpiF90Kycc4QXwL1VrisNx1R0Zx5j9q05IYatHg
+CPBi2A65lmT9dH8qRlEvPofg1rg3V42sqteGqyTMfa2xgGBI8l3MGXeqvsGQaE2
R4aD9TleYcnUfg3/cpL8ET1MARehxG1jkrlnU3nlPIIrUsMk387lWbUiI+gkHatP
KFlMaufGMhZklsipKacY5YPr3E0RlxrfEfuxFxAnerzky8pe7w3l70seXpmx5jsB
v8eNmMuUcpRyppHXBWysfXhNl1AfCMYp21RLAEqvsZYt3/BJ5gfutBup06qHsLZi
Xz4sYu5O3Cm7pXUaxq70am4JlExaRXZwIidnjTVh14QrB0W7SQ+Aupxmu8WgbY58
1JIXLg6vHVkLkoDjwOcbDsPnhWSjPoxpesvidcNUTtI03TcCSWoKDPqVS2FCTjgv
POh0nouKjQvYTfZAtgvA3VSDdXTrPow104WuRG6dU4VXQi75g8vFby0ci7q10VBg
WI8w50fuXlhkYoLsaDrB5ivhKrW3RRyYN9W7sp+/mHTvpzWxzjiJeymrMSC9CgFc
UbKzPuXzTecer/XblSDKeUmUzKga6RgfzhvgqCbDu+nFl5T4WY2elvVtT8s5V2N5
+zv1sPpA31aTurQ6Hm8bpuc8mwUaAbJZ+oy7BHZMwSGibeglQ1lpKrSmtdsGIvr2
ysxiycpVmL8kypv8OibNIoJubxBkZ8VEmbvH0QghclKGGTPitwsAt5W3pc5r6Q5W
0FlHRNg7Krw3i7/clLGn6aGeyeczVWE3GYX4FzticStag5WsLxTY2viUWiHV4FAd
tCMdggQZBb4wc102EiQF6kXxrEiApFeLvcc5590+npKU+DgKkb2vY5HcgQnDk0h5
UkWaLlWzi7E/gto2w0Rt8FWgrVMOx5q1oP/XIgIUWXZKqqwxuIVrouw2467tUHIP
HKM9RAK5n/DFA0RoHWNssCZIEwIJoamTTUzWQl2M21+7WzGuaNcZJ13sxoYT0iUY
QjX7RG8nwkqxxf1tu0sLFJZWJaNNiEIXTq3tnlrQ4MGdJlvE8sSX6zQBq8vaHmAo
gLTVoJFb24KL1U83r/k0OBRb9GsI3h3bhAc1apA92UY2DXTUhi4N9aVwH/VSW53v
0dfkmUGm1yAKFgaCM17DnsCJG2vKdXsQWnjhV0XiS7IcRBj3AC3Xj1SzM9MVTxsn
OYgv67gxkcCtVQ7Ezt0nejUbKaXlVzCo0WzU3jWwHCEgEnafWJxt6pGdcOsa5b9m
GiAm+Fh0sby+SxNNZLYkrVklkQBdcj5SWJqlOy+wnisgtzXa2CL14GX59XEDvw7f
BUystFfqcruo+PsB6ZYf+G2qA/g7+WfLhsp3Q2DX7x7X2/lb7HAtBhEQTLjwmxj7
ubYWf3OuaOMHchc0fI6oaJpmmFaEZ+cbz8qA/5qDiVEnTLrwkVPRL0kqOEqvK6Sb
itETR6KFveqadxxfAMsT6zJ/C0Jdxf4JEsQuRCNDymMvtGVjk9EXDEsEQOsJ5CCN
Zx39d5V/py/2QIa9vud6ucLtPk+T6eQOlb7KUph2q+63yFitPtf5C/OAVt3M+lrM
9hw13LLWwBZMtNLVy/OjdcJuq6XQDNn2ehON8XCP6DuYVjon62BogESYzuT4UIV2
tCww8trEFmGnOGfqNSB8s20v4ce65SG9RveENMJeG+nhLKn9XMWSBfDd6Ov3emNc
PFAl7mgRKxAuCWRutnQ8JKPmITlkITz1RCeNyg3YU3Oe4eWum04sHWy+d/0p2q2S
V5LtkpdfEWbReze3jZlYW1mu/aFNfxInnxgaKWLwKRdehxWh81SHKKgCnA2bwV5H
ZWGw7T+T6pNnvlCKEnNX4k3yAeyGoyS78igaMb1Zvyz2uvrcmNbXTTGuxNfh8b12
0VeGdm0OEdZXOZFFBKbbSnN75SaKg0ZuGvcIjW4uChAxH8PooMnqYYilMate0GOR
LBPYs1t+fZ1acRyISrF7bPYtYyqBlnYJMDK7SBOlR3sl7nHWaK8a8xkWEuqtifJi
qM7bwgJVDeVYMT4D1O4oclY6N/ZKGVDNoywKh+4kcijMTZ0iyK1HiILYMKAVVhfw
vC9Qzr5ew9GGIm/9Pjm+hPnPQWyoZMfd4DOMwzs5IdJi0cEPMHaPq60uYWBp1YCb
pWz8thQ2JiCS09r7+/sup9qyYdLo9BMYdGQaQibuphmjkAJzq2bLjaRVINaPNMFV
dMfVkJBuRrwjwEDJXOoppQbmAgxfNB+uhdZn3iIQv6gVfveCIzWVPhZ9tB0XD5Qn
9RNb+FHt74YFzSDv2VESTQZtJLcU0QEw/Jf5+/ydl3zncAYlKzlcDviEfkOuzeib
cFPnm3Mz27a3yorhoHQAxtOtbINvqbgHoSc84m5AKX/7uDGV390QOOMy681JGeWe
ds0D1QBZ6K2Oa2l/6IrnHuDQ3YCLcFQ8VbUa3AtYrHUNLnh/ynnKxyyiSm/0vv2k
syKy2ZglKXXRbnmn9eUsXdMsEEmgfJ1EDY41Bx9cSiHABPaAK/JmpLZPN6UUxTz0
qupyEXZ1q4JV+an21FoAVjPwipinkK+RoFCYw5juigrieTd0HKxH0/tq5Z7OW5TY
2fuAluZ/UAp+zRtJ3+TRXSsoCHEyW8Bc7SgJuH2FG0/tEYI39QFukI6R5U2SSXaK
x1nfdMauKrmgoOr59Az3kXBWh2gNej947r8s39JaPhZRXUffL2zHkqnnrcOAsKzI
+3PWZnrRR8kV2qd54zRVHkFQwpKFAEm0AMAts+GEsw/VZd7yAv9awgINcFeSTmg5
YRqt15k5wmTigTf+BnVTRZSgAPSsxdCnk0rwdX6xFHl17cMKwH3pU+wijW2rhsg5
6TTJM6qpRyxihOK8JzTpgvkEd83sH7eK+1BKNlS2Bl2pMt3yvX943qIFgsbLP3e+
OL30d29sNMopkTwc62t9YOwbkfJIRykaOYWbPdRuLvh3Meve8gIl9R/O4rXHDuRm
xyCqprGTAE2F+btt2Bc/LC+7TLADGW36qgEBfxzGw10e0DTYBrkRoeAGC0POIhbe
1UFwbEyk9+GbHoDWzGT2SQG0erUXk/krYdmtfPKT5Yj+SSdzjs01+/7qZIDUcwWq
DvMgmFlZPKOTxowG95tWRWFOyMiFutuC0NEzMRGqYTpp1S1Ykw2ZQjywfToFqUFP
nO4S7j2j9qOhxCzHq+2FH5lhAHDnZSOskyc2PJCwWKGSUWhOXEQmnnjnLipYA3gs
W3lvIUiVSBHO7prbOLcqIqtKm/XKAhePjp6MYCf2YZc0pnY67D+laiTiF+ni9O9Y
ObTpNVb+z/qtRq0q3aYLeqjz45QuEOkGTxEL3rPGtB6i2b4/+APUvvbI/MqZqJNd
YbeFhnqPA2LQIuJBFBJ4rkRqinkQ5hu6RpB0+j+kPOKGjY31slekgZGmvCgrYgTq
bHtJrZZ69b/Zx2uDjuv8i6BmYqHSPPsLYAbd6Ebt+/qUeKzGeicHsN7tCne4lpSk
wYe9YiJEK6M8LOlM0cQUOXExeYUUGMHR8XpDHSbxd7zi5jnez0SFbeOKzG/iyiMC
Vml/OYBrbFZ4+pqJP6ZYzp0vyKX2jSuUPAGNqbpDDvTVYGepEbNrVew33nKgDwvP
w/zDcmlOZa8CKprjbjrPsrcBd06pYXs+uqFIG5shBevqbIls5XIAa8WeplElUVWU
YmM/76zm5HqT0t1rBSbgJYvVQbnQF3XDGB0P1sOD5OYSgRxXgUIPxwqlSrVUfCAM
D0uOTT+X7KN/dcq+fM/jhf45HjeRyv6XFcdORK7FKsYnj9f8+pAwK5wen/zDbmRw
lDuxvbNDpfW8uYeeLaX68PVDkNNK7xylTCIUaCjWwCSeC1+OLKRZ094yB9elcON9
yBqssx85t/L12CiBwGDCXCCAduOptwkfXFMpAv6ehgLfRb5OmvnbH/vHfGM9vmHQ
1PLdy34hWEoRNeNX71ZjcwpK3HgpUlcNW0F2of32CYUy0BY1jJHV9MTiPeE4LJHI
09oCr9kZy+AAvmSw1xPbs7d2SDPX+YAHykbFMyONYfNV8dTTOB5qR7dYljDNyCMB
NdHjnGm/U41WPsYMGwbK0P2mfjDVlYf5W25r0nqdCQCOhhCVvE1GUHbP9Rc6K4jm
2fCkZl9Bccbz4GalSYh97IdhdnPX/EX1hqlDbQtFFpWl1gcddc8dkwX2NKXcv8ki
BQZ8INXGP8fJ99pe9+a15VMxNszvhTljn9+F7MRE9GyYKquzJunXPHoT0RAh54HE
k2MkRdmyqGxvAU3qN3Jbt51SG6cu3BzSImeXDIyG8wjUZnDGaTO6osGvdMfKW3Eh
ZvOobRiln+uBmb67bZcwOKy+ESNxRazFoyG9WVslse/3VkOdzdwrbzps5e/GIf/5
TlaLFIzokJedGbYgSrOo17jLoFVloCa+Q4DnHveiJo90OFt3oX/kPkltIcnxPRT6
S3N787ZOdO4zwjgXJOEDpnLntBMrTTjq6rLKFQQE3GipMmdvscpKQIFSzH9btCPZ
6FWitTg1JN2j4JlQpCwUZzxb4J3sq9Kojw3RjD1QvXAFp1Giumh8iMYeQippRnVe
m0Vl1/dSqmrC0f6UwkDlbEjN8lBesIWkcQ0C/+L3wHorqOC9PB15ao0wS6wZqm2L
SvnpHx0sT7Cs3Tcx53wfDIZjmZn/6bFFmpm6fXnE89ZFE9svcHUgFVne3bv5t/VZ
AOFECPscxg/0lhAJZPzaDWdKOnrS/lvsPsuQ44LdBL0XourqZuP68th9ewW/ZYni
YVMroPbFHzH1+V8x3X4+Js4dlzfgyHFMfmgKRsfGZxQh8a6sTSzt2TBck6ePd/kj
qRG//hSi13wmgOg+4wZpuYu/FI29RPpV/T/NmiM2m2ZrnzHXusvZdKQaDuICbMCK
jBwD0shw47qn4gUlOzYCHwlmJj7R4u9J1XPMvG5LR1tgnOZdPMdsCSzO3rFos5cD
MLMC81hefYYjxQ8xqLxArpG/6LLbsqTE2QbBRi0qk4I+QwDFF7TWgEy5Dg00iSDU
FVnP+tcls0j78pJsSle9tUMPOuNqtBdZKlRoB3McJyJsNQKH2j/5aHs711K4hc83
c1EoaPpFuRin7ORCewSTvtwpYkhh09dMluJnwpCS5dKkeuPgbdDgM+16y3er9x1b
CRGFmEnVlegg+JGCOD6IjkiqYUAYpuEcrniAixYqk/6Kbmxm6vh1BUo09W7euzKD
q/B2LQPx2fXGdJevA4FrbWgdaGtspkOkpapQh2oADcOPr8rDLHuSOU1T9qxpUtJ3
YOto5revqsbkAfurMer8bAJkPkLRijfEPPWVhCIcjfRvZ6aysrV/UOoW1d6dCpIV
I93g+aUTkZ+adOtsTu+kQ6yVhuifmQUhQEJJNMmxhGT9SlQhYNK1oHuQ+1pVQxgN
NatSxC3361uM/+sY5OopxiJdAuPpwGgMp25rSKnyJpGkI8RVZmRVQP/b0WZ8qFuE
5YIwYFBaGb3GsWAJhwQkbHmXz2sVR5JkWw813MESuTb+Mva3nvy3DGPlUAboK+rR
SgEDZOFY7DZImiKSXSRzLsfvweqEMA2fOOcm0nn25cL0pvwA8BztbIC/SKs10EVm
T9aTkL8v5E4nrVP9ah6q3iayQtCmMmskFtPnwleT/ZH1VGq/aKb8Q+uKugmNjpUD
yDhE/jMueVSw/5FRRbj0ShPokv4uLnvuXY/p/K9tFV49aMfJwKYs0NXxDXC38Ll5
jkZgQBbP96xEL6Gw/pxjcmM2CwnjKX9l/KQ0OAAYZ4N5UBfCMPGDa0+eapBA5xqb
PlGbTUS3cOZLWebEg1ymIZt53PxsUJcYb6a9niXqHDAYhxHnax9vxYlEdShqOp4z
tQgQVtj3im6xw85m5LeEaWD6cfdxmWzZBDPQD6tJDKJeYafqed7gpviyu2UEKX9t
YhBC4UbAQMq/sislZfnG4A7H6NIR3Awuo/eGbZmRJF2qEgg6optIpvmFcDRpoufa
do96jVpEqJdUuHUekZCW/FDmy4IunZNVuC4LEX03St8QuUXT43d0Hy5cRwk2TwOQ
fOftRHN7jOFRoEvFeQEdO1C84qAAjJ1guW+EZ7QW/GIRzsmZ0EkUKhSdsNBpeY8P
GJD7+QaO+Xj0egSIeSAmTPtUNqToEMnfBkID+BIDbaYqs08X6LS8ivpObste60Zc
c+9fLcryGbXVA2jKKArbakkAroXXYjn/zfYozq3/tSZrd3lVH0dgb7aSGdVtgfpS
d41Y4r+zNT62p6P9P+DbySnWVap6NIrKUyScC1JitQhfWgjjNqOO6n9ksBOjK/b5
q7wWckP24HhNKTOhh6ZqyfTOXlGvVJFgdDIjMI7xbMeIKHA4XVJDUZeEfobDTkp+
k2dTdVHMgWCnjbLwre7m3WkKSeJ9ebgXq45B81IlR7SPHzHdDq+xsv59IYD5QMD7
UK+Np/PoiqqIc+X01sptzva0Y/dQabgMSzVNFDAOY+ZzmNZKOp972aQv7YIGFtiY
/aOtr228Kjy4WilyH8bM9brNE+KEgZLpxLbMflVuKMEOGT7gUx6AS7HO/Y3rLKxY
A8VMrTcE6iQgEXhJWet49cRNo8Wf30sbOoK1vrCdWDJIl3bQoSqOfKruZiTyaGOL
gFYxgKgs2H2qeUScw1s+nHOBNvJznvbJf3R3Tfd7lYUWqtQrbzmn+PMmqaU2FjG9
dTbNQPxtHwT+U4rHQYO4kPiUFbBFPSqQwVrXQxpgDGbb3kwCdt+VD5sFZHSurxGk
JcjLF3TpXw3alzXr7OknsTOjGXDelpjk9hc/p1i2kBAfCiZWx9c+3Nnb6Xz0A4g9
xp5QdDlEG7PzPMzVzpG487rLdO3f4QsVUXlR7zx9mPmKsuUOiFgndDJCiFpJ6FQl
AI1y1KU/4lE1IYDQqNPskvX/MK+hzQqNIBznw7BriETnKwarPl4vhRy2AW0eCYNg
5a6cFTYzeRzjBifhBlT6xVfScMmMoXCOfNhuVxS0Toq8NuLU9RwjLrDO+JoX2xjm
Uj8FlyuMaQ44daNCEyPJRIUO4QMZDtynme00AXJX7r/Q7yzTqH/xFt5ODHssG0dE
BWJdt5pLhy3AqFCG+z2t8AReQdK3MUpTBuNZcXxwoEWg/marbGFDnFOUH1gMWm9+
Eextb+TGOLIpvQvhR4rYYRcfVcLOZcuxn2mTzQwXL9QYhFuRzG+HutlxQJXcsL4C
l1J9oDaG6G4Lxn/kQATjsgwPV11An5vpfF0R2Z85JftDui4ewODfFSWkGz8N6ZWj
5invt6APlCsbwWP+P8+helYYV6liyhHOiTUvHQOk/23MEQ4ZFSQdrsxg11HDdCuA
HHD1+XAIPZmcs5ThuiY1PGhpCP+c8N5UHynZHvOWKYAltFq69sgJuTaYlNk9zqCf
D7T5uTgp+3gYH54CP2Immn24Z092HFUQLdDoGvSavKRU5jgNXdnrtPt+pubFVYds
KKiaojISzggXkWO+XNGNGDWHdNuSKcn21VFg66QSJqfPG1KD6eREbNOwm5fEZgVI
JnK49ihJE4uNdTbayhsLUDwL2lyoITYTauc371CY8hZUI9bs9ZgY8VPeTp9Mkm2T
UTvLbNDNJZ9gfLtAK9EPebezFb9BdhfWPy3CYKB81BzPCZUOXBk7Nssi8+CqZzEL
zz3dPZQid5grxbc1+RV1DcnCZZPtbS7CGQtlizyuAUgTnMOIYqSBaebrZkyR2zN+
isjSkgMpMHnvNHZuW/sAARzkWZawKn1Qhhk/xtoUtUN2KjZMLxadKaDSal/1oXhH
5lWgJjP+wE1zfXSoK5fD9GybxE6L4+3P6e4OJLy7qmfyFz/Q9ue7UcWKLKuIO2He
LcK7oFNMf+wh35F/L+3QcX3UEMoo3hmJgf9bIzP922tEy+YvQchIuBrCAnNpqrqP
OlxrxTd6jFqTakJC04b3/FzfpjP2CKfqsuzGyGGmKCIxfNu1UxH1FHDKWD4yfU5w
cUBuMgcvxDvTVdK0JrouAaJtiolue/0TVplxp++eqjso2dqE/XdlBun1v5PSwZ5Z
NaTxusQyYZYJ76SyQr7z3+3fO+InvbrI9WJdBAakZMQiDWmocbhjjnfmSOnhy5Fp
XKq18nDd8boaEsmolb6L/2oGXHNqILGN1YHDQ9xX0A1wxlrq5FpLm9d5DSFkk1O0
IWKwFwR8x8JpPo+d1wOz5zgREyebCdaJpi88uAYAfS/xMuxVT5YrcqyXKreiUkL2
9DxBgsTNcL4AbqCNysNXLz2jexusLRTo7IICSe2b7F4Xypd9X2Vwigm9MgR6SudS
4BvQIGJYNvybONo4KNIOi/Yzd841ldQGYQ639EWV0p7vuxCo7qRbcc2jqy1ELmQv
p8xNiveEI9FWjPDPLQMDgy0+RLfpeNRZGonPQGwaAKkSR5y/dCE4rr+zsZAUQ0gB
xAWh7fYlgHNsOuTy+WUHFNO0S6vx8eMl1Nz6ZtOoPXU9wZb2QHlbKMo+ubkmBwk4
Tqb7cZaoht2FrQdzcKsjjRgmGEL+MXPLPldEotYyJnRu53Nr1LFhTJGcVbvooPTo
8vAp/Nht6tblzD0tW1zssTKVakrwrph47P2st16LrLpq56UWXAlFcSwVbolhmyQ6
J74TsJKLjAT/uYf8a4AyW8QrlR+XLsXYK/9m0qhRvJXj85OcJebVC3fmiPEZA1U3
hdFUUmTc9WYo2bykT3Z8V7gfOAjtpMV5/gZKizOeFsCHDKscCcSSTopPNS5Twiq5
kGywG15/Dbecx947lvIUvak2/UEJy763GmjJwuk8h2NjMgYbjc9S7porF9EbTQ3X
QMVcZuDZnfYJ1ixEwv/hXTjStwZ16DNHOPDVYKflf5UORP/dhvG2bdtm3nevL54G
XB6QMnk34olfWRyYsZFLlZ4PlRM7dxLwZMT3uWF4vlubEXSz0hYxiySdwTugxhCP
xwI2XQCag/O2Ysb+Wn/K/+xSQBK7KbTdfricEiMAb+YwzhyYQDQIeMm7bgK7y/mK
Cf9AsMPtZel0ptkk79e0HFKZSIKDt5lHoGDik1YDgkz8BYfuGT1ROb7wP3tlByf2
xcv+aYz00UETHDGHjA0GhLWerbFeyC6UF7Q7uVtDrbIIV4xHAkxBDkvhvKe3nFZy
YPQIRwTrh57YBpDy94wWjLOgPds69iKU8zJOGShUPnxgWMEePglWuvfqOY/zFiiS
5ZD7gg39hakyCfKMjh8ytHBR3Upt7OmN+k2KOauV7hVm1BQ0WetXTnxsp7p9SbI2
d/WNx8vthzEwPUxT5gRb7l14Nufqr4URYhqElGVPyZvQil42H6wXP+A09/B0fBf7
r/HO7ifKCCXdcpFqhRd1YHvb/kUqtyNmWCu5BlNXW8qRQrq8XkxlGjiBtaipZQeC
gnsmYDtGY94P0yX2sFNcKFjoK1z0ZmM/yaax6D1xrJVZX7gJ/sOBbkQuQkDD3zp+
2FOZYl/50Mx3pWNK3j/PoO7l+zny0Z3DNAHPyuzRQGVGo3NXuOqXKmJiFuWOvecG
hIONtxAzn7Auvak9TeBO0xcgGSaiY/8dR5FqEyJjbSXb71Rzho5A6NMuDTRIkBiL
OLUtedoIJd9jFljZmR3xCZXloHgQHKDx+TNb/9tJNuFJuYVFT9LnZKiq1MpEutyb
Vp9HxVAjHUQinTtE+HEJFAFmv/X4DLJRSYcOYPg+J5dYBpS+QNTsLP2ycOctWwhi
BRkuGfic5Q4a8fLyY3eb7aexWgab5TqL7zhR+0C7bKbpTSApOQw3cvgbRXatPUXZ
gniXjUzliVyk83NumDWaxuCyaSok024cC+dmtFRCOw0cWdLKKfYiZJZ1qC9McuMY
GF/86ik3WmM5Af9pVvcCXyDGXcmRCYQgwCfrBuSHD03jUwjU4faKWbaGLLEnO08A
eQDqGybxXU8iFhLCwggDDWvWoQgGGDt2o5dID0WdUy/pZVCzd6SyUvExJxJlEDr0
SNWl8WR72OUXTYH1Uc7SlqJajOiwiPlWymbnwLPP2+6WZTKKPmlkZvLTIyuADtSB
b5A5/0V8Froctr+VrG6hZQAA2F1uczZubVIufbAYIYar+h8aHuFuUKUJWk7kQrRa
E8kQJ+4ig4FaXuxZL/gO8NvkQJDp/OAC1qZHzcGOVg4iDyFVHf0TEG0ygglfrZ2H
OLovjKxfVTEuzPB41ao0Z7LhLPM280cLSAdd97UtYr6kcO0C3FCE0uqHcaWVnUuf
zoQnG4lP7DV1W8VKzwvKqeFNtOM9L1n0ZDe29QIS1ADR/ZmaLDoFtm6wrgZXIWSZ
lM8bwIJSUCdhde6EDzhiHnmzLPPtH7B9ifJ1r5Q9hjdur3AJtLtXAdkVlRbBslyj
KAo6ngfj01+qxBtjbz0hlgvsgJhH1jPea/tzUGdTEGCpzLqO7WOoidUJtBhjC1et
ToxV1me04Exc7vonD4vCcQwu+X9hstG+l5BxZy5OL1HjGKZ//5XpJY1unjTokpjc
PW064gr0GW/8kAhCwvmbd/xYz0+AQ1EqkMeE6HSeXvaUf3OhUXnsT4ddqI6poHUy
oh24+lsG2dA8A5MODb5rmOrsOEhzTJTlVaeY/fJ/qpgI8iiJ129TL/uLMmL7/aJM
IbnH4gwSPE10dVYQQR1hLzAQSPPMyLmYkKhh7XtLOfEeGrlx+EJNXHbhboeMed+8
PZmBmlFA3Z5WXgZds7lppNM56dCXp+I7cnV/3X0C2Akm04xtnU6V8WsOIbl2NxPD
7f8sK6ZUYhhdghpWZZGGEVHjfOeTaTUQUsRefuPbFJjXXLsO9PE4HgleSfd+9kDV
+EmO8Tcr4ZBI/UfrAucnPNIRb5OqoMyJ1qD2tAKetD4ZQIsRs2o/NcVIOGnpBVkG
S6yFGxttT+vwNcohgRHGv8e/uJ4E+U4MtqWgyasMBI4i7iOK9ekAhpsbAnLAVygh
NGqvb0Er2a/RV/vPxzgioHG4VrRwhuHoRWA77F5PC2Ru/X1OveTf/oLT5sMKMBuC
p/2nciKMD2/vHmI+4gk+OirEcGbhSyqTyHNgeYfXgh8HXlUuUEnn1y+aJvk6PGkY
NMyUKvQ6PgLR7f0BXl/G4HYndkso6znpJGqNifeALYOMp26JaIG1Y9w+GZCPSSnZ
QQP0XMS8woQV4XzJyavv18I1HAXiQzcq9Rca9UEMMAs+KE6L2kZAUb9Q2OgNq6JG
k1scB/6vX1/s7T7we52rOH5Lz0b5Wx6OxsrZm0Uxi2dMIq6wc7icHPXwrlTJziL0
cfqyjnuOU49ZQpCtYzU2q1VbAGcpwsbjnEX3B3QKKdZaTc7RXREu5NUsa8cZTzzA
hnm4ht3qZogRxrStQjKhRx3u4vRL7xCnx2owjMJbKy7W02h+Lbeh4w5gWVRmX6Wd
qI6RaTEc7tkoCyMMnyI9PRcPkfh2Pb0tvDLxMVOUhJLf0GidyruN5gATN12dluEF
3OtcP16vPAsG3Ikxk3kBzZPE6/HvUw2oLRHJaZqSEULDVzl/IbnowyVThtuGverg
Lzb1MHv+v2W2xRcO9RJ+5KUZHYP8DQ5DjBh9yfWIBwseelrTBJGzjNHIIztCl/+T
DCAWDcDkDYscaQAPwigcA0OZUZEkcAExrDKiX5qz2PCXhrf9MPmzDGvK1HBtB+nY
VwR0beDHB8bLaiOizgwSBpk+fkNmqcjiqWHzkQveCne069w2+Tz0MO1NblTR0mSO
lk8w01JNIkiTyI1tqmqlQ79E3ytv5Jqa9d3AQpWwNCu4yz9p12UJZhrsAtVzow66
NmBuYjM6dpiwyhTSGxLU8Ok9uTAr4znF00IFhQ3/ux37BprvmVMlRf2G++SIMtV8
UdAjmWuFJxALVxVfDt3aWmO1gQ50+idRKPg9Ksaq9IeZJaMHugTtDllxQhu4Rn0Q
EAcZbIO8wui0U1GMYR4N37FcJIISNXnCKQTSp6+gsvcpptHPHXP4By+3gZ0HR7nY
/LWjnojDK98W7Yn6mpdfcOKrApW1kDiLhqQCDxR1bFf7SPMEjlZZKJ+38F+u/ou/
rn6MlnnnGqmG1oIlEVHr+hj4wwiP2K9M7uxq8BvZ1gJj2nlYfvgdlaEsQkqAFgM4
CXO+EkqbOJWsf7HZm+qGjt/tyRkDOQUKegBBPZ9KVti7wNIR0W3bXtRYAdBBuoGu
LUGLulmNXDLBLukVmIX81z0tJ47NCw+w6ylwNhtYaojmH8jIJAKKapMRPmbWm+i3
rwmIHzDG+cXBEp0FHPlYiDFU1Y+3v+nnE1Y5DB1mA2BFrV+uH95TDcB5m22VZHrx
E4GknarH1w2Qrt3Qykl8VWLHAd0g0BOOPpkWHSUWY8TpDs2RdE0BqALEFYCHmMBn
w7nfLbJirAXZE1tjLU8EmgkDG+vWraRQcCItNTfIUKq5T/pY9AfWVS77kHCVj3uH
csTYthREzPgKidqjTZwAHUqm05AGX9mtLqLn1mULxMuQVXQuFxDo9iktCxe90/BY
iMCYtoX9oSiKPpq4wdCxU4fMoUH6HYf50SVPDrrgcMRFw+7+PzQgq+sI3po3bicr
v6lpYplbaj2Kqd9D1UcIyctEY+dU4jqcG5Vj+X+aUG6T2m/ugjr7ZGlFQy4gxSXu
K0O2Ba9eR3KeT4YF4LmLO4KtBzFRJsRLYmmrc1oVIZBZX3vYRTklDalj5d8UzXrE
Gms2Hlyafwfcf9DI1dUigUh32wgGJ72uwBobc0r2BsTYmx8win9tnMk1WCmAm6ry
9hj2RtBTKKj9gJwpB2l9VhvahJi5wwIC+JZivk9Y9r8CUWhcRNKJGcjtQ99/57Kd
BhIpmNzMOPPD/HQeBINb1sY87qRsxDAmdXfjDkJPQa37VW+g3UuCPzEWxbkCKqlB
s8J7cF1TcKEDx0VGXqKxJzoTaYifId4kmi5WysIIGpoNOYcoS5dObANoOZ2fLoP4
wvLw1uHWbvGr8GFlerkOWV+EPvNJTmXJgsmJ3HNpmtvV2LvJ499N7n2kjN5BmX/V
oTqkZzkUo6lhY407RqEFSYd7WKYKn1eoEv0OIFex4kRzTkF5yrKUrj64cOteyEsr
M2FueYbWCh+ndxMlgweNSd8sdbIdX1LNW05Ozdv0z6XX+yMq7mstfo4aYF0lMDvu
8yHmqikAQZguo1neRT/YKkx1HRNVx73i2UxIYjnsO2ldgVdPf3JlPb5MeL0JkRDM
DBlhbloNEuMCJxJNKXybtQ7gENuT1rmREhzqs0+/MKZqJ/V7K0nGU9TbV32Ls21l
NeCGkir7XJ3WrWVbBK2nMfWrGshzJtS0zs7mXVbWuZyNOhSyr6aX6SIjNV/IwVuv
oJfX/SAPyVsNHHIShCO5st5mqMT/55ZmTHcj5cRvTu6kFh9HvBT2hGZSl7jAnKmS
Qphi0Lma0YFCQU26uFNBz434q1glMSRUfFuWkmImCwVj2Ru+Bo4LUzUHJHOXdOke
4cbcPP8ZkgBBfAl4laFXHLVg2TodzXVkSxhQIlLyxHuwPK8tG78uzesDz55nNQsm
ZY6zdOeJnugkNjS+Bdt4SA7m9rZAACxMbodskJKCBQbt5CeRGkrPnIVWfQi1nOZn
/leodVj4vyNyXDx3A5w8ccrTz8XhX3/pRcwU3VtnG2Q9O0EZP8aQ4Sewov/siZuP
dEx9Ef1BlaA8UKRjmMkBXH8dJjvpLCus8fzmxHYftvAHTxzoxZAk0FvKEKM6aQtc
6+njb1vKUTGd8ffvNO2pCtD43FIgbtdtfaIx8wKBpLXI6owE7vGHvHf96frXnFsH
L392XpXwoAXi1wdEfqfRbx92+1AqrRqnkhpVN7sqO+/3MtSMIXuWLKDSoRMhSLZF
2AIE/iDNeqhAVs/6sQaDAaEtt2HROEr3Gw62WekDcnTcANxFA7fZ524QTydfAKCt
bZVJ96UtKiwxLpX6R7FQTd8bTWlF662aMkW2QhTqWLfAOaPZ2UWJnhpKHM8JyCUq
fcfOX2+31SiJ2Tg5D7qh2/H2lbtIb2+2AxWmd/bjnCRM5bDcETH/jAF9PyIGj2bP
6MzYyDvR9G/Gll+d47MmR+oWrfwojLFoxOQL+DxtNZxCuEoLVDlyoMIAvsgTwM+8
DF1Q8++N0qDuCAgP/ECOM2K+HeL8lN37duVmB2eaG+zcSfJ9f3Fp8R5tgX6rFQEo
X9KELLtZb3yQ3SiLsaBxRVU1PqB2rme/HZuGAZ3d5HDgS757wifTfa2uK1rdpcns
HvmCGPgzsRkT3UQ31Z/41vSTT3BoOrPNO2ZcV9U2CMcPfc2THhXZGeKGQ8sZ6dco
Wj44dCqz7k2wFP7Cs1BO3gyNp0jTUpCNpkJJ/v56HEpMS3ao5LRW/tC+g0siCebY
63+wovpb7qZZJXzNyT5geNwl4EiOPDEIkZo83+8Z7QQmitHUG4W2Ub2rl3Ae6buu
H0gF6tVfFcBYvWdfRkndpcHSrhGjjBXAWAcJUOfbV+HuEu+DNEVIe8zWve6C46hm
HXVdcYiT4xhYCAZC8vN0MweBS4x5DxPurDs9nvn6obxp2HiZAHY4Op8TU2zDT16B
+kPfGW/9kPbamd4PPUKM/tWd9BNjpRn8/IIAfzdXzjGxZPq8v3ks6e3EyxNVRWCM
e10vM1WemJJf8yQBu++budZpDduv3Izt6KEznQ7f/3ovF5qShrHsDAtLOS29VKql
UMa+hg6Se9r1UYp5rRZuFCz7b9JFIamxRDH/ZSOPLDbBrQeaftpnETZSi/PDnm5j
s0txUR6JaLK5E387ojrnmtW+jqunXOb4DtxHiCFDLX85Lgw16rpMscmEesNMKHgZ
zMgH+2IG23iTm9fMSXEejpWdQCdnOJlC/rJ9VKyScb+TPe5I+9HYgR+Io9bWFWMt
GQMXQSAxL7lOYYK43l4Umj7MP/FHcVriMCGqbK+UabHS0ru7MllmGGh50IGvGOPh
S0nLcgOCM4h+jC4lZV+O9TqKsP5UfGwCwkEu5AZN79I1xT85+CXFD0J21qQV76cb
PV3kyiBuPb95ZGoIxEMj9vjxYzRYqgZ15SfOJZpbj0gEjG8BVZ0lFR+blV9vUrW5
9zli3tv8OzFl/pu0n4iWY/VwQ0FIV/upvjFBfsxNpgp688LAts2/2m5bsfEpYl9S
mrwG1964g+kVkif2SHh12qtfnErr2lgjFe7qpXRnNhSCaaIMIjuzvH1vccl5rNEu
iSFmdTnoRaZDmJSvdyFAQd/ti16uOUNw9tMRnkvhlkehZa/tRb4VF49UACw62pSf
SpFKN8Q9K93QXabFe9QlsXYTybjIhem2CjdcDunJJ9RKw5e/ak5x/Z3G8KDYgbck
5JalAHDCQ63cACuRLlGgw6hWkdhN8P+RKLBaeDQErGCMgacgp449IO0xKcIhLNpa
3OeiYuPWejUP9Sng/+dfbKWm1GZu9nvPN8aTUkodsgOWrPfvMaqbE28CVhTcxiWL
r1iPeYghz5nATRfJzjkURVgyuRYE2nIcclvMBCIZDPzIX80WdYUNkIpoQRXXNvMl
H7Wb0pK0HAxxGXocwDra5dk0j2dmPP899BjAPokZqOMhfyzEleJp1amAjMbrSnAy
PIWOwjKW1mWr62SP5KGKhS79ahMLcPsfE/1plodnQ1on+3Hnikeh224L+zDD42oC
EChH4/Sj+W3Rcm4YBtwMHKkgtM/TVkfghsKdA3HSv5sCOlR7s/XT2A/wOOeaJbFi
RpblSh6CARhG46Si7tlPFjcRn7+5xczaddYAGWSOEgj8jMT9whCzPiuUswBzzFbO
yvpGevTPFCk8MW+YA4hPE4oscSiHCi53Hh6Ae962835Vl0wNpWZ3xPXytT6OikMW
9oc/fSKzYUcZw51NVo1xMvqZQRBAJ76BFZ8tyDxm2O8RecCsUvkh2zYNPTwFUAUH
AYCRWcOQJlMySjO2ikR0bse1CCTiWMjEZhNfdCpbg5TMpkmADiQUaDpPt72kU0eL
y0M/5hmDqdk13T+SSRzc1mH30zV5LVaRQvMlGbFkIs/7kHT+X/r0KaT+zByPHUGE
+BYWJKDHAMRz1YiyHaAnzw5CYLcd1wU8GBXQ/i69RwIaf8n5ERoSTUy4smYgj70i
S5F7AAeC3n6hvy4r/fsoAoLSER5HvSMP0kcMbrW3str3Za1NGLvar6xTdyDbkptg
ygjjJ40+k3NJ1ggtv8Mtx4KP3Lj7u8xpqLnxjr/e8W/g5SIS54RpJovMMeuYf9zh
M36PqaOgnfSUU+UvlPqUZj3WmZ+utWfa+bK7qq/MARz65W6PcRldhJb8sAiYBGZM
HFnFUGwVMA8lun8aUi6J1UodfoVTFXabFAT5cnR2122LBuwtUpcly5yGpVOLKtvi
uujfnuiw0PUhxZx/310tnUUDwMydEKDIhbSjH5Ci7x8+cKKA/QuL0Ks1pDV0aIj1
B1pDSEuujyh6Z3yBxv8aevo6yxRFK4t+7dtt+8cEJdWs51tiY5fUhtkyhjTYFpwI
rbcU2/+jtbVk9Bbnix9ILmfGcd0TV7EDKBfSrI7qsqyEY3VxWzKY8SqpP3UeUzAu
/uRU/2QKybSDDYgXIKyYsEbZtCGe43imezELzDZ9+Q1nSWd93kr/Im8VpHF7Z6lG
+a/BKGRfePRbsWW42eaAiIPsdxrcDQB8pALNEI960BmpFIszxla5R5mwHsybuHWx
8VMLQBdofg3pz80fU+MSmqTNLJG4zmdDgyf4a3U5PkJWiih8C9au6s52y6CXdbrM
urdkceQli76Wkzf1SgRbLlN5foZBde6/SeN7xuEMJaBIes8nH2GyiTcS9bVW+FNo
xWuwP8wl8yNI5b68RsF6Q0qNKvcE7n7tp4w/WPOu5xTuInZCaET0pfkh8cCGQGxk
+xOXdlAAY9K5SAqBq6IHL8ibjQL4U+5gimlvo/DcKCdI24U9xchYKWH8bksVcfDJ
zy9F6IjxSZf6w1zuI6ASmJqf4rEjRxQRuraioNL8v8F+Zr9wKy/i+crn5MOVbkK0
TOngducvCAGHcegTEKmJv3C/89qSMg1+ZtWF1X+5D449kUSiMS/uxOtUFxicOhk+
Bbp1FcYxC2p4A8nF8645DgTl7ya9bk3CAHBMIthsf2AqPiMKYDGw/Ba/aRq6S0J2
OwKnzxOtoHOuQsu1bBdRLK0eUolB2zzMzoKOJ7XAX8D2HDLIEzzNNjyGaZ+BO2k6
05wn7ew8w/e65HxjjM/ke1KKvMPuCsrXFgfCgcefeNEKKc7h3D5F54IPtiY9UtGs
eYbaM+znL2LmlgzjB+YZ/976NTs5wR/P4wkKvlD26unCWCyQPbzJi+WMYbSHvL95
snu5hS+6sUF7BoiqKoMVJE1Yu97C3kZj10c4YJGuMmCf5zBDSPbXxipOVbyhbOni
rA92RXQmFQFIab7OxqPjBUKJvoNNK4erlMJUDm2u7byD7wi9qez/bvlyOU5I946s
S3Rvl4I9EWb865PxpC2WKRMlgzR2WDBsNnQ0I3MJlhD/REFcZehkmUu0dWd6rsd5
ogNsTWo3loVVt3h+ifR7H90Ck+JoeEFbGPOTxCnqvHhIwgM2+oFLNfmQPQIL6EUZ
RCx2Z4EEGWayYVSsUimjuaDBh274tANt+3GGRRA6/FmSHDCQhinxrc329Ln1tNZ3
5S0LzRm+l3TvwbrTM4x6rodCcV+XCXGoqQtYcM5n/HgvHmdD3deAWU0WfSUT0eVw
BOt1Zc3eDvlxwx8OzhMVTEwf3G7abcwI1v2cxpSRC+M8PUdxRkKb7p/NdD0PKjPE
Adk1PjWGfFTNJukXypfKIydzQK99cozTB2wLwtMb+cpei7l5eiAx1CRhu5PAD+4E
0uj3++aD/9yt8910oWly1eLx9ZI9fNNsje5hVzo7DXmqjukGp6Ys8n+CFZGiY06U
xxjgjn9l2Nhtl8jqfMCdaAdj3wDA7rVOO8OSGJqMh9sdwW3/qV7ULoCZ2xynlitB
5KXiORhno903qm6yzTEWJsRsGE7AFSakWsHXf1ey0DwxrGoBf2N38JXItkD0mc2k
SgfoEita8v053SDIBv5viSQLLPBbnqI8xgUoMhShmnvltmWr9od5yOtH/lmIzfyM
fr2p7SjkJtLGky9VodwPwfCuQa71SgOon+UD1ZKavVqZkSunTpeILx0iRV/sSDq7
mByjmVCbIYdcUh9doCtywvwtoMMgB9Sza5ngUUZBdXI+aIbGpJxdfCNjCJgnZ+yb
MtjJjikr+phVsVma/w2j+emGSzOvZbHRxw5VK4+XHSB57O+DhbrmJEIODzHOztf6
5dZQprmc/KJH3ItKcfSMnsyp8eZs7pZPVoOdupvCc2iayiGRNaFsllf/Se6fXdzh
2i1sLANRyja5Hw0Gckv5xzSxUbEFTmGa+RJ4owYYzNM1Zz4MG6GIH5BM3S2aGUZy
sRam2OgmuQSH2zPnTxkHkoXLVw3nJWRimUssxZODlCl6xwKwc8RtErGKzHLtQ/Gb
KuEKlgSOdG2NYbx9tGFPgElhFJDKqr6H1i5qG6WxKfmcze4f+bu4E30/lRX3YcwN
gJ8WkayVwV85rpn2LawwoGPB75H80qvI145AUMc0QwG979COasvkt1mJ2oOV3jJy
6A/RKI+YN1VkJ4fj6+sPicJRfl8SzHP4vQg3AFtkyIqQMG8vKjH2ot7VivwjvwkM
GE0AbN08dTa7ryw6+LFP7wFaI1d1GcjbID4NuXziQ7s15UsShfX9b9kgyDsMo/uN
nJ/6IDZ0XMUMB7GJRJppknupuFP4I74KXwiu8sTTECYwmUZS5ns+rx0iymvFHTBN
A5J34kWKUWRc3F3qSimk44M9sLe9TqbQdIFRwWjo+R9o6+sOcps+Lx5IOzdHLRW3
70L4ESpj+RBW3Lqxm1oXn705Volt2VRpdJj4YIliZQEprBNwYHB6+SY0EspdhC0u
pPQho71V1LQ5cnHdtfnqWkyU/PfgfWWAUwwIseYI6Agb/mhhfgSAq8G9cqMWmss4
vA0dM7fYH5vxa/DkCyH9hbi5GetMU8feRfC0tK2KE0fCO8eruRdbCInGWdXIPkWf
6hWHXDLQ8qC6+Do0CM+TFXaQK07Ls1ZeFvm5ISjL0MOnR0z/Sft1385Q+VreYIQv
prEG143P7fd684f4yEaR/PGGjuPPX8nCCIR0l6iKZ+Rg9//IwsISVQ3I6g/XtPDt
Un1Sr/7kXjRjRrQsQ+mXVbo2iT72nJhILn5AaJOQM3WYfl+cPpharAkJdCVYkeUc
6x6Q7kT8Q+a8L6KmdHVaPmansg8Um9rRctePjSqk6yp6tKfqlb1Ry6A9DoS4Su/y
qxWFeUsNNdGsBF08ybIm4ro8jPOxUpY4Nd4HyLGyFtioJxxU3TR+kDxiHyjroCNk
blyjLo+Vocz69hY/eu0ocRsAv/vVV83aoofg1RuJoKwGhJ7wOxHR5yc1nsmeFCcU
vnwgm0tIi+Q4XUt0wu9QWVfC0xazBNeKYND2NB/lyeD8Mnf99SSqCuFTJ2dp9hr5
yWtQvL0ADhHBRG+LTq3FKvrjfHOhcbpOenE740kWDGNmHed3WAVbqVYj3HnnPP2/
R7gU49D7cB/ROc3eMaUOQpAl5IusRPu2JAfoZTJErRqOyKTP4gsZgZZxHVRPZADn
3wPYgIuNY5a6M0Das6QCUACKiSL18IoDKmiUSwkXIRV/blBWVlTFH4cB95xJ5YAu
vA0TJ98FgZvmCP41P7tAyXo5oRHEhDDNnqy87S+EvVBV3SjBAvFzljI1VeLEX8hj
q5uARx6a4lFff12OoFcBCdwang+uWsEPqUh6bPcrc98+3DtuklWXQwgnatTbwAmd
kAnSxJgxWe/ytPRmWH2CjR99NNDDjnsXB4EkjoQHzs89W+8EcL6Vq44m9ecgt3mL
FP7+7OyiLlt4ZScA2d9Hxjasa65qC894sx/NClMOS/BDkwdaD9RBbAaU5BULvele
90iVliR6pJIvVPHhtt4hpsMCLX15bwjk349BOVb4+WvNosLmmFFfKKvRsASfXuix
dFYkhCKRp8otHvXb/CJcMX2zOw9GSP0XOkF28FSbIh8NcGP1Ig5RpU+UZKWOJE5m
OOC4DcM/Wg/0eiNswA/1LvbmtDzkyLgpG/Iv+uTtdo3RiUh349Fqnd1TMt2FXqTo
Hyis1W2LSD3aKwXjklh4SjRvf+aTbSN/h0TRkcyRRVuAp2ug6QWY9Z2N8R9kUAGK
K2BXskOFS3dtnJ7QgMb/lbXMHSvjD9TxbjjJOt8DEIRseWwxaGn8UD8vFpIHvHaZ
PebLnh8sLYMzKY3vFc8V7QbmPE+DCU3vsRpC5DqbP0lWSovp/kC53Ad5B+gz66OA
P7OAV4MA5DCOuYX6dpIRfJi3y6tj61sHi61iF4PsAolpHuuHWfMIK5Lx1ROlsw99
u1wONIA2snnIktEhTego21QEqbr2VefQgSsJAGSbI2TpS6LcBEoMg5Q1ikY2SBY3
G/Qbw45qNI4vJdu7LPZQpNrMkr4AfIfAd0sUGkWzvsGrZzCwCSGCh7VIpkYERstC
e/nzHXYicJFx6Ww9guSxPtldI2Cb4n3fz8XGZzxuwG6MJ+2xaYxj8kSDV0xWrY57
gPXVvX9HQQCem1PynbjCqqNiCGFxqvYUXIP8+NCgNrShOOtyrKIRYDHxj+95zG+9
CKhiRfsTkXRcGFLkmLIibB2uUUshraCj1PKBVsnhekcXBQKsb5D0uSff8X+eAR4r
lc2ywhF2uMTIfhpb35dI1eIyoGzQ8BYUh2nfW8SOqwVdWVQ3EHsOg56nspchaLVd
KaobV/mB6Q1b/Ez/RbB51NZbJsUWIDzIBZtSi9CjsAd+hlZC6Qm5s4aP9WgL0/p3
YA116WyDzI4B/s2pDuKwfGPXMwrMjO8nADsCRGpYXcGTahrfE27c75s5irwhi/Yv
QITkaplU4VoNHFtlWZSsNoqnNLpKoOF5wiuRKVBa3s5Tye1ZVw09xDVeYOfx17ba
sCbWmokXK/bU6Hr0XzBhEFxMjavLqqDgbL/EPUfRATvuKb7A8Ld83eKNekXlJ7XK
lh2unjDASkX8EDBSp7jVwQzJDUGDgeUSGozSARwfmTD21g6A2vAYB1PB9jP445hO
UiYBT8xIiQGK2u/h3zNykx974VcogNO7ZLcSGb78lVlLePEkUDuxia7HB0I1fuQR
GQ/W9g5cegZM3UVUMRgNVKT1SzFvvcTxB8yhiS0xKKqGaqLIqjiNDYL3I+ekiSID
+mVv26r/ZtiK4FnwPVoPYd7Snv72nwKtVZGLpHVkrFz0q20q94xFaeFjNqNY3QLI
IlV/3Rt2nh3PoqWtDYdeDg2Ie17SioMx4mVr+4dwfRnrLhae6kgaoBxP7RhHZI0K
Nddw+GTI5HB//ABjLtZau4DOD5qWw/TWUsc1J1HNkoaUaNpKjLkPdrvqlpePJyX8
BIheTkKdOShlzke24a0THwRj5jWtaf6UihGyF9CEJ7LmWj69BW52mR9PMGklPqa9
7mXq6Glyg7/nkO+Hgznb312FYjSCN8kF7ydQi3x8pwl1zPmePU6/ojMJCp03cZ0L
7vsuv4rAC/HEM8UgCQ0TqEjpxdjoznY9Djk1lgDFwx8zlbW3AAhHhZmOUoNYBQnt
65dZ4M0tfGV+VJDywGFakW+opW/plDmWyae7xds+7NrcWlge9Mf6TaYx4Pboi88i
N0YQl36Q70VAwk6Ir9GKwIZEvw+a8UrlrEZHv78mwStmggQsHmRhf9MRsjxWVuNE
sxgIxhLojLKs1fdZrao293lL6mEniejEPO8zwUNMveGFg9WG/y8hRRNRmQPgLPOb
KAsnHGu0atNOb2b4pW5o7bJeMnAvM6Yv9tN4KvnKe5eokCTAS1wx4AdvRx3yuuZ1
BBZDmsW4qzC7IoGy7emEm7RzdxfK/TzdFNGHfRXl1lEvRZcaylYhucRFJvQ6xmwi
jQ9JdxauTZdqevkXmPVEsFq67FfVIaHImwIW7o1Qt/FClfAeY74zzigeSOoBlWJa
GHUW0rTIlMV1iNWFsNhofZvIcicWrhOI44XjNwm5wjVJBHa8/oLBRj65GIHc/UNT
sFRLdiFDzhRFv6Yv7AEnfjJlboycTq0a/9kgO/dxMc/XbOoOh2y2QI6H8Z8mdGWw
dJr4rPC/33euC7bMhTNiuSbvNCf7BEALr9wLXQMkerFIJgnTyONmmpYCc2qyhDJy
Dvx5Dl9pqKzrfBhyj9fRANO5OJINuWN+NY5OKzZR5QYHkzQ3Y+LKxyRm/wUdENBy
QLrgrbJd3B4Rg+QqcwlFdonNIdpDt++X4aENMq/p7jnsck9mfqCOGsqEZuzY8PSm
Gqbia9GcARZO5XhkE/GKmmOHvHVNTXi0hRg+b7ixx++khM+nTefsB6Z1OFvlNu9m
SqtJjqbfJZ9TlDXeF7AGKHCKUrCwvVNWxFg2cSPqf26nhk8kv0+hLeI3564F8XW5
BNCZ5T8bzDCQ5InDGeSLTfyoU29awOnHs3LxjS68aUUGECEnSrhp2wKqPLlzPRKG
KSO5OURqEseHERtmBXJo2dbjY/o20/FjnsghKYPHM02rmqVHjIphExIORxWYboKW
oDNbnBCabqc8oAUJ+iaMmcnju4jpnUhQjqBnO+QNuXdWHtJb3oV7YaEcEtGuIgSW
ONYhVDlJkwdmE0CznuPrCkEVGqqMhz5i3ek6GIRZRvVDaaHsjo2hfZLabjWcdUMu
JKmvOsKEa+s+xYJPXIKJFMsSn0poJzmyN9mVqGq8oU+zAgwhs8jBeEQjHRHOHNS0
Mefk0NiJCrYQYvzE0Jl5o7fIEmFoJKavRGUgDEugVGLWKfxX/Gus1/Iszvc/rF3m
s7WEVJkzrWdsIzVoNRREgXvGA7PQCDGtQIGeb/MWvGokc51c5BqXkD3VaEKgOBBd
kWV9SjB9DALWfASD3uGgp7NJ/buPRGUnOXEgdOGMfwb4dfMdlosbrQ8U7TNi1aSm
7yDZ7VSdPG77GOf7Y5aNmFM0TJJlh5Oe7JiAqdJqHk/Z20gL8jKXeNb/RGvp5YJI
IWMuYhAcPwh5QB6pgkclvOgdLmpXGlJ+HJEmYSBtWG8wNs3WA4iYhsOOTQ8fslto
xeSBXBt394v6mzuABEjZ9jLjJ2yAoT0f7sff/PwCm2FFEa39ERfL5WCBQTUA3Yzx
i9ilgC9SOf7mLsd9vyfjX4+RsMIgBWO+sv7lnm0Zn/Hzjg/G1K6cyNxsEEHskE7A
s6uYRyZcMKb/dF+jqGXlnc1TceufP3DFHazC/mVEdWGy7fAC40p014GcamYrp4+b
zx01q9tb9NpY5adlofqzyP+u/E2mZ9dmIB6mU2MHdNectNZoABWkzafSqEDw5U6I
ngKtn82yIp4s27Be2lx1g8HM1+pqH37TcWTv76LS9vjA8fPRDMn/32Vp5HtWN/jn
u+3Wknn5S63LSHQR0DTXAbX8GMGHL3wfUap5oP/4rUc3MYKephyAXYrpxr2QoIPU
DGYokH61y6ovBi0eoN3z3rMCMS3FcR+o1x0uY8O7/SUKkiMInXgva4JKJX+xUWxJ
vhlRBuBygAH/sVTV4ddGIyUzXYBGZsAs9LND1/AdRgnJ6J0kZhZd4yimhNyMAlSk
kU+I1MGjVpDCQeWcJPd2Hq1MseFMCzH9/KTnWsye3LHVX1QsjZtvfUIgZDcQWWRG
flpJo978vqrA25r5iH9UwugM25/kLZrOxg+C53k84F48rbZWMLAnR5FNhpKWnIzR
fkqPLNN/jhClwYDujMPiml32T+36xAHez3ly9FRv4fIwdSzb/zSD4O46lBq74APc
x/dgGLIBGjju/9ZDuh0GVO6BwhuHl9DmfPGSM3wS9ZrewGQOqLNpy2/Vdbcx5Fko
+dsYlYLag+wHZSsoGf5BCuHPAX5Qrl+dmUEhDOAaPRI0FLpEda7+nL2bQY+pOdRv
53P8p2bUoFrjFDZxKz69RvohT1GtAwpJLfR2s2Id9wSW6Hcjqp8bKs0Fxi0C/W65
83+CmvjoozQH+dqsjYGwSkGjVPQSxp5T1P9gNmvhMz+fGfrdLbJry1ybpI6qD+SA
ltZGt9++VOncQ+j5QVK6lIwnmXuY4O9YuLZPZcjRhytza+6su+iH0j/s0buwnmxb
tmLzc3x7VI5zQMbyRyhkn5S+ZIsR8FzunzewFgbdE/hr7Aj2E5FLxDwuw8MY8wWo
gFXt/pTkL/jQN4atMEIb5e0HT6gJuaqWx/a1dB9Gaqbi5pjAJH3/VmTeDpGWyyI+
gCfrPfL7UrOeJwmX0XH3/SA4Wzm3lSfHP1HQv6TFgfmWR7NFLABebfNcHK1Sx8y+
s7YIV2IXPTuQNk+8ANhoihwsCOxS4sQUcG87iIaPagtsn8D5fQ599W/3FL9vCkwi
Ip2eST+tg0086Dc2bJRx5Pp2mdjEOEuT3moz0pgxsJg46Cs2MAwLS1Wm9iCG/dLh
v+bsK0EeQ4yxdJtuQC/pin+rKLkHd1VuFioxJBPBgacJ+wqL9r5Jn5Gfs2VntI6w
kagywFqX4PyewMv0VaTUGBKirZ3BjSSgx2eCxXaVop31JLtrHSc1H2n9AxTtjdr4
IsePv5rm02p1/3wSDtpkBk/Sedo1SeC608Q8gC8MgbG+/8995gdh7lTQ+O98Frjt
bPqzMtKhqgmjbZyI+Xc6iIBhs77NLV+uSp2TqV//66JKo6eSMZCvfbdJiKTeR9ls
dJnHH6pEwG9zL5Q/nYRN/QpO7/t3s2ZOXI2VDhRKijYYvctF2Pt6Tnln+AXyd/hm
TYcKMXr5MBd/2TT8qCBfVxjpw0AGA8BEriGjo+qD53nzw7x5eXL1Cksl3m1qipW1
pkDDs9bQ47NnSUVm+WQhNf/1h5TAnh2MZj/6aAYHSgcbMH9Zz//taHkyaxXYIovS
uiyb0Pw3O+8SsLVtvPJLQiSXTXQMwjv6W1hj5GN6zWAT+mhpZzn3lfU5NOU8zVoJ
3D3Z/dJsML7nxjSYj0IpEErPYnP2/v1yGOXGSOYseV1hwv9XkYGtiYZvoWuDcIEi
i6jt623m5+ZPyU+pegIN1levuwh6wkuVnvmQmD8msFl3fc/qS/IU+rwqXYFABXcs
UWqEchYK9lrQZTv+bVUcG2JAzio5x/3q0yM/Dkz82ePLx+C6tifdUQNyeGoZN6/u
2Xb8s1uKjiO4ckfJDNobetrL+TD2Hd+4AcsAMaphaXOwMNVhutywdAUxh+pCghH1
Q1BADs7DMzk9Vw4jXjtAO4oARoFfGKvGDhoRMN4K+0xQCumqHXxPsDyvMXlE72b4
lHqahlLo0fD2l5yLR+qC0QJjMcaMalmYEsNmQkkLOgwceaRZjkMpnH3mh1LrWWXL
QhS7GACN5CltQVrecHhkhgKlPVM8SyvxRFl/N4roOJzNm4C/f7YD+BDDtA5t0EAF
V8LrtUOz94ODd/qD4kcKLb++2OIbfwnoQlRmLPxYR0zYDpPGq0sa9/h1YimjSTFs
TbM/rfyZR1cERa7nWgJv4T+QImYoeUYmR/FbIN07uVxdFLVfh9RynAxNxyqtXDan
+JP8YGxII7jTQY+hsd2YKCHwVVYe9gpxXF+JAdNeb/9X5F6SJepWUNblGhEzbtZy
qFdfAJzXpdOBWIkn2gQss01HR4JJg1/dk5KFa+jvdUcfkZ+iI5gAJwV5YONorNlT
ojtJIDR2ZSb0mAPe4VGFx3FYDRI6B41uh7+our4B6UGo4HXO8pplQ27i3QE8lBli
XhyGsQ4TvqrvsyP2tozZo48RHfFuPGXxU2MFe4SYJ2BhoqbvMAQ9TKOjRKgoAcU7
UeDMVODgNUQjb/cdGAnbzokyTdyGejSfx93va1V5+JCo4+/3x89jJq1UwcQBZRzs
ASLpvwcJMN6hvAen91Zqk+0UDl8eLva/+Hg/cEQZkyQeEQ9Wib0osFz5/t4sCAhV
4AlrqOWXZYKM6tFJqSGHvAiU6GJ3int92aeqXmD6lgL1ShfhIanMgxLJW+ag3PNv
42x23wXIdp9r680s6nftUJwc+S8OvE56glYZ1cM7xY3wALOINuPZMR+yV6OVV6nY
DFzqOTyCnfAdcJQATi5ZGUNIFCBG+oy2V0GovI02QYAGH3eyXmZmD3J+q/PY6pJ8
SSfG1fBYmOAxQvbj/jFYCSD9wz6wVd3QXHyprWvAYMdh3JKtpkmzNizhcC+sHXD/
hrKX/KHXGwDzEfEr/1sGWbo3HiqVDl2uHNqAv0qGN5NGChASULybf9MD9tDTsJNX
to8aQron8/MqTKIztyrHNi+7GySwi6D4a6TfyaPo5xSjJpXKESWe27WJ6xvE59fE
KElGS2fkyetag8dKkAHqxEtmr5wYQTBaco+ilbk3kMd1PjznjTZSUkheRz9Sw0hR
hn6R3zchRByH/jXzodJ4E7VQEmOmXfiwjyiYXi16ULLmffxXN3ronKBdZKXglIqx
0OOSkjQofc1aa/Weh6ozd7ovzZG4aO58UR2E/nWIug88H+6rnZc8S+8cqXRHOWZW
Tm2ZV4yOuY7PXahFlZngNgHJTbxqXs0jQabD49KMhnNyBs1LmUmGMOvPx+rgZdu6
T5mw1M9tjaj2oy1aWHlsm0tfQhAcOv1nb+q2VJkOSyhTr7zUa7Ng4m6Hv/XPfxfw
F+jJ3Cdb/eVtbiK63fpInReZvAv0duUFIds4c+iOLk32m1lXV59QjhNBM0xTSIpf
c0lRR81W3bU8lrFM7u1zaNFicp0jId4PCpcBsB+HL9aHdltXkSBQRSrDhY8ApiMV
LuEPoTZPELgcLDjdEdo3J56Oj/aRXOAiyx1/7E6wV0qQzEt6BzQX9xQrfR2Algi9
ZN9XyeNQ6WukqaUAx+Rw8y/VCtN/0DJy+vvCxLUER+wAr6ow3Ih8zyNwGD9lShwn
I7by7ypp8U+NtfgtYE9W4wnFK9J4R9/wybz2Q4Js0xlDR4Kixs7H17Gt86FyPW9Y
Vk9D7DXUXR3UiMAW8yFnlQ9DK+fGVYjkpQPKL7tIz2/DcEazieCRf6np2n8Aluww
hP9UOqobfNd964afN6KectwPG4Gv0bDm86jbN0aHiX4bzjht/+BV1dHCal3zc57f
26JfuW6fhBGI41boLeTeb6u8J5YIN+AM9IJYE87Ad5glMsietJAV0DnS9AeTJE/G
iifZ7OQPPMKNGI+xdR4aFPFglFt9mmNBhSd1rwcxWZzDzq91aTUg5dl90Px73/+I
nE2xIZUiBoRuPAKZk6BzlXXQK0AWLCslH4dlXmeKRUhwLAuu/230lklVulu/psK7
zpnUZ86psAHoDTsCGzCSN0JgEi/AAJwIyTXDQS3qW0jiYrm1QGY0QJcaaL3UKRwc
O8Mf3U8w1tPhdO1UgscrTV9oid5oJs4Wa0vH8hOu6xOuqW43fjBCL+4ah8D97lyt
WiIF00MKY1JKW2OkcPZqlRdQz9Ev/fplOKoFM3Dh8dNAzSyhkuL6zI140S81sDkQ
95pnqzJhc/xblDbJ/gls88b4fgk/kKKV7BfIYdniAd0GzUA9J16pDOyZII2ZRRQJ
WqND4yb1apiWjYIm/UPiwTxOG9C8YI/O/QBdqO8WYzvMmjXl9TjxyZNsNUbVaOzz
SSd0/jDDe5WmmOvuM678YQMRZ/OudHH+Cx45lWxAdUrZmbKsDg7A6zoA1duKR+2s
hZlBATo/KvxCo9DniQWLBTXza4N5zUAZ3ZYZX0PjAHc38GXkGPhwkX6rfBCNUCJ+
zQ+6x45sWq+C23wKHU/1bgFUzYXE7T61mTODoqOi5o//UXb3RGiV9sj7lPBv5vke
LH/MSQBcIXr6i+sogWzkAZf7E1bnTjZpVOdMQ6U4G5sKL+1abqScQXNK4Ci/odhB
hH6jJXLDYzat4liJ3/1OmYnh/jEmOhwCWC/kJ7MdaEv2KWA4PJt1p0EoPtGpwUES
hWJOnfuEWnJ5yAx14jvEEIZjS4/AjdazYhsU6QVMXCnWCkpOfy5II+U4YaztHBae
G8CRaaFeTfZg3+AONrVZpGRylwrftYpXm1BGbAfmUX3sZGNTZIEXCkCxk8G2F5BZ
zZHxZ4Si3snJvWf4Sk2XAGKVkv3QHkedGDQlu/vGzi/ni2ZvEwm3ICuIksGn1Smp
VVl4atfyf9k3mzyxQTZOQd6UiX2SPn7UIdYhkNhsuotHQ2b7hd7BTv6wxZ4y/e+a
ApfRC7ZZjhwSxjVTI9MzEpgcgOtdm+4lTt03EjDku0RqDDqMy/zJ+YHSn9YyhggV
V4w3fM7kH235W2rQ5Ik6NfwJ7V+T3j7IJx6i7qtd8oHtjFSrllFnpWy0HvNpKUXl
s2vPI+Ez3yP9TTtKrQwzjQPJmhNe9pUC0lF4GRQZiwuk7usVj0O2VIZEncvQT/5x
AQfU3mRPkAvD7PExWNacmyGfcL3WWzuZAZMAoIgukqEG1NRE2f013pnKf2P2j/lC
4Ah6rGoOWr49v3vzo7duLL//2PM4XMwB89fpeil31+cexCZTAVTzdoZH0Xb5t2tu
yhMRhwCT1bkGc5aJqB4mtz2GfsrQsBh8QxAsK00y5Aw+R6X1oCfSUX53xy9E64Dq
HXo3Pj0viGxItBsDDJLADTArmlrVGbyseDD28pxDQLmvntTCMCkQx1+3xoN/WQrR
Eieksq2w01KUC5bgEuc4gY8AjvbnXPtWbrjZcQvubBlnLLgdtM7OYFp/2Me82ASw
ZuYDtgSZOt8xUTLtQG2rRqk+aj9feqbPgMK/Wzprw4aCs6Rb6/c4IJcDRwnLkDBQ
xbHC/0XaMtqnLhhre+OlbMnEqK5mTPk/gYs5py9A2D8riBQ7mt1ct8O7CS/wLt2Y
0PbILofD0UydrL7EAMQ0uYSm5BMdAA5/pDKDFzCgfM14LNe2JcL5+opXp6MUOG1k
brtebE64hNs5gYKUNTy4CL3DGR2fHwCUFMh6aNGgzDis55PLlsW7zU8mw5T7Qs6L
X+96R9nCh7bScpeGTikD3/5BBXPJucYcuS/0msklBwEKwRrElksYJeNaxjpzGjwv
FVJ3B21sgJofO23epdTWt+ZaLx2BqiK0U0MeCfMVwpERUi+RsEiNIOY1dwSFSWOj
KdJxI7fIwijQ3B7+Aa5w+SqHOOcC12J3ydSOcMFi2YNod4OLUOYnpdWRK82yP+PN
vfZYnke2eZ+cF1+5TpGCItSJAMXSAN+1Op9My3fQzIUqPQfr1JXEeVbHQfn1BSmP
9u7btjK1VI7Xd82Z6eKHS+5E1EBcqYc9R1DAzYe4O68+ITSD/ba4CTKBJ2319scV
ZGbvcf1Bbgua/U0K4sN/7GsnDOHfUXg6eUXV9ySaH3IdaC1sd/4+tcoQzSU5NQvK
7/SNtRNWn7nvs9tVpIQUvHpOlq9vO9DLYrtYF/JlQiok66I70iLYG3omn4ryudzp
6C0ixCot+Uh50JKOE8oYYPfV/ngutJ1TLXZ/K1nis37kUnkijkHqoWHuxRsGmUBb
dp3fKheExeRP+B+VDKUlqCeazlw8UriRmQ3wQkBv3sNerm8opqCRICDjo82aQm2X
JhotxTRLMgcz/kwKV/CqrEHYUgqvonixhKvUk0o6Z6Om8i1aljGtMNIAw/5NUniF
Due4KcqVePvgBSiVAPFZVa117Kgw8Zg20nGFeI/kluoH25KZF15xM1RXm1awXJIm
E8spzxWeIwDYuy6g0iTtVGp2HKN+AUTOIf/MugD3xmcEnoM7qsTKlq09VGUQ0QrO
89itM34KbrxbouaKuRyUm856540LfUzItRE3qyZzzYMPrus4GzkqizvN4yVMXVow
D6hYF+9llWagHvsKmr4REqGWKH1A/V+LbzDdiOcpjXX8y8YO9ZcvXiYgWYHCIUHF
gdDaKEInAyc9d5iXLqkQH4l2GQetKd8ZE1vvEzVmc0JRyKFR0XUWb9wSctvK0Wa3
16FykzDXuNdwvKxbA6NQCyy4jkdO0V5yu8YawG8Gy3OH6JApPGHntcf+0tTyqTEu
Kr7zkG8RV/EddVFnkBXVZ7PGXdYdCn0y9HyfAPMZLDT1PUheT9dhgFOWYLOuyB4i
tcuPH0wvyiDcr3l646yEAUfJdC89hWcsFbqnBVN3MULkgVB8hXr3mMONwZidPR5v
FTK6GTJYc8KPXSfvImQJH2Jm09RCB306m9k0WIBANbepQNOBcQbt+uyeZx0RZkdq
gvu6wVmt4mEGfFi6IhB5Ol2WLZMPRVbHNLf6NkIuCUjWy7PgKiu+e0LK2cXC1bUx
sqXGhYsm4IQmarScZ9zMZCRnjoByzITAKHOmdpGQc77T2HkBi2hsFP9xxlNnBlpI
AWIUXfMe4ip20maD6ThorD+A8RdICZ7MfCCm+Sw5+WCswz8ERC0eUUNcGI/4BxZ+
hhtQIJtXifpkJsyMWJlKVr1wCDrub0O0mGzMglC7N+asA1WfmT02hDCO5npIplDa
KT82NxjwxQjR97h3OaKrCWd+W6vev6O4KuUys/XVWT4xoY+jRvyUVMqhUsX+g2Ub
Aka4ceUKm8wCYhirHX4jYgI+vLJyWYmQPrgKJI5a0lO2G/udWtjgXt3oPWbr1gn5
gZ/eGbDvZgKjavicOJO4RzCBQATw0FjxKaTl7KLmm/IBQ2DxSX84pmqQBxcywJ1K
ngB62lCepa10V+gr/gJ7yvpxRUdDluxZqKemaZ5K8XvjQnosjAi8UERkTgXQ5y1t
R2tYkSyM6AVkIp9kmYryVmk+GRtkLBvsWzfe/ieX+2ygMKFCE+gPYfoF2lpADFKZ
3CkD1B6oGeyJIyjU2pjJkOkMNO0t+U1pXlYnuek5hoUAiw514pRYoZ61e88ixYCX
y8St95EPyU6k7QFvwaIdca8JVQNmz6O1ynoar8aZUkmAfx2DwtDtmn9a0rqswH+d
BgnqVGyl2JLyZtiYQvvUwNS6UbGO4ggsZFe4ZAR9vuOmIhFGrhpXEtnWPfDRvLf3
+NAE8hnaT9jyK4tEDfRt44OG3yPlk4uHeeMumy6pZgDK9JKHEXHzJH6BXh3D2oyI
ZtxIoN7frufvN4HGUKvRqwKuWyYTHRYe8ZJIv2dSgPH10Nm/B8eD5e5sCyCUuFrK
tfzgI5vSaRv2ET73c6+uKFu4PvcpuQT+P1PXMxoYu7y1gmbWm6yCDtzBEtq/b/CG
QDagaqIpAIbUPgh//XFKgosEO47L6gEh3qq7gTd+TN/WjLZck4BYybTArzHoKZUV
UuFTCbr/oKoKLBpfxlkhMoJcU7CpO1IVjhkDVlet7c725fLGhFgT5ynX1OD3O57O
b57cSHiN9FMVVMMN49jpDiyt2tLPqgwag3DQHBwGFWyEpLHn79wEH5Vg2gErADtE
oxNf5PC5Y9j/OqwpssYYANEd6PB7KX13mQyBBogXC2PWuNR95OshBr2FUH6bV7cj
xxzqQeE5c8tumINKhEnhxd5evAMo/OpOA6vQ3gC8uYZDxzvH8T7eXnj3ox06KmaQ
+QFzhGSv0wg28TwKF9Xmg9iY2v4ztmc95oa/ZdtGcIYMnbt09WJdOd3/eZwLCjAj
6Oxxv44hF4ILn0Pi5evVrVYJqjuCk+b9s1LuvSLKmWAPCIYszwEitc8LNyB58ei7
IFby6TDTtFDVJ7kW3Qgo4lP0XJLkkI6zjMrP7Idfiei7vm20GEb7RR5yif5tAV3V
tWJqU788v3C/qw3P0l9d9iwMQQMHNl6iskqxjDOO+G/7v2/De4ifTQR2+buOGL/5
ekwc1y8fAAv97n4BxyH42TONNNoV8Sc52HRGv9jenVSejvwlAih/4v+s6Pz0W9b6
URvSKzK0CNGKmSryQoNRdlY/m5NWvKCrtTiz6ndb5UqRpsMk+2Y9sublnURlWTQR
WVt4dA064H9A8ZjfOROXP7/PURuzFB7W/wL9ywSX3CJ0HIq8UsNSW7wphiVloQlV
LKSYThgUIvHgWVGVoE0EIv2RXSdI6AfKUVbogi/8w8JCqZf+h+x7t5jyxT1bzYQO
79zQHlM1x/ZQJYr40oTs/Q5kqdbyi9p6eOelT7FhxUbVojh8ljlq7mL9AwHH6u5C
hwkVtCb9FrC8n03ExPTOVECZ3/E3Mf+SIQycN4Mol2+mbG2TZcyuzZTC2f3jfAsn
2tvxq6D28LHkDi5rtJTHpqeAHEmguIj4UW5HD6F4GQVq7As5h/BUcbDRdDH9mSxz
HIc+aXtLSvM3q5yI5H+9dR2j/LS35fpIybfYVehled6DwmrS4zHnhgSrIg/+tGW2
1U+9/pFu05LKjjCAhje0dHz1AyK43e/0GrAPIWqTn9489tKLQoHo9Euw5B+5CphJ
LRFtAz5g1kU/48Z3B0pt6p4Mmu4GTpf2BUIapDGIP7zy+Pcy4pY+WxijKFuF/RBc
yvmwtLLsonJJXnE0fat0gXM79pwbpfmtMpJVxnwEgzLP5D0yzX2xQwk5A5kRFiJi
k80L4vuKNumV1i1Anyq8+GyuGCQmY/XxcEaN5PWuOcXumhbj8D5j3acatEFn2/QZ
dPfIZHkPc1xaaTUeqJIVfB2M7nJTt5tLVEBGg3v5/nvrSVDQAkJ7oL3h9H1wNu5/
FrH4BemMb1NPP/tIwtbIPZMQsVrf+RpuSJ9JUfzIvpZgtloRhVVWGdncOL4/gl00
PlPlb+PJVdsfrHflOwIN1BUhhZIdnswtSAn8zObjNF3/ESMmt2D48QTlcLobk/i8
0Ewy9boGev+/j5HXyfU5rjePjIXfQcvSYITGB54jREYU+tNzvgvvT/nvd/4fiQ3v
dwsnS8TIhpjeymdDU76pUwhqmx0qH1b5MMGnVMEaZ9KFZe8L8f4LpP0+Fgg4D66D
o7Ug+QtWeeQDaOPxPin00mH0tDPlssTEn0J+cKS8y26IWiYHQTJYj23Ji87idC9o
R5vX/bmD/N1dMi/+y4MWKxVVS0sHjlvJtHUGUgltRhoY0Ojyh/haWIHHR/0g47qF
w3/7SS8/+KnEa+N5ZKCg91DNFnX8MTQRggaqw0Ml3ur2bbEoMx/BgHdMMqU45k0z
tZ4qVsEzK2BaijorKUEcQtAchUCu5bWn4N2Jov3denp77ct8Ve+rqM8V2N0mduev
ij1wFwSWHccQgIDmXF5itr9DOq07XkFA8STAE+Xd5iNZ40DyUnuU/rA4IN10nZam
47DXdK9HDEgpgwBHjP/sp1FXmnQ78hbmXi5XYiN3h57bDSqtY7LAJyXeL0XyxH9Z
Xq1FAinhnUPqFJ6AHXCodABWUm47xuuV/auqdYsrx24RZBn+uDDpXi1liyKSvKuJ
hnFW+y1mQvF9tqNyDiJiwWG3kLtq2QfS7zHBIVbCNhJx1lV7br8Zqml78pNdBunt
McDjtLwVJdaK7a3lL+iAkdPLNTgd1pDi4vL5g9abQcHBVXq7owN2EbBiTemU3x/g
80DpUmKo6K1kAq508zH4R0cuYZb1uWy8aTYjHoni3GjoFZK/xRO+EwmJb9ebHeUx
uBwGo12DjEcRvVvjljKO0t0uUoP9HXQ1y3DHhkF1twDiUNI1WERDA3g4NcreCO6n
tkZIM4e7urS1+dSjhHt9OdXhp5AnMq5lO6+NzbFSn1rb6Ov4qx4ZnIcmA/PRy+++
u7m/2SuVK3iGDszCnuMp5IemVuj5OpfVeCt0UhWrs+fJBe/ihvM3luIFuPBkt9PH
Bv7sihb42ndjS1Vc+zBkrkrnCBTeelfodg/FUtSY/o4+RPV7YV9KBi7uout16/Pq
Zc2A9JUWynrqBtO+KVqjdE/9WmU8zerWnsdH+MH5ocvRXNDK/GKu2c0UjcnHqMzA
uOidZ53gbMaSVXPhMbQwi5oEo1e9SHqmVKmNKmM5YQW2+Tvv5u1PiehrhjKo+BUb
WczEAGYDoI6EteeYAyWv3cCVsTlhUF5rxl4HZSmXwckmC7E06sM+ojXgsGfmmH7I
E6G3oaL95et1PJcwbnbdtR2m5fJR3IgY2/78GbG7fKKk1qoKLrIzRZn1At7GyXcG
icmR7XKSBzHBsWW8LHli7bHdjDbEew7hXNQLb25wFW7vzSYc0u5Za+k+nutb39KC
R2QtzoQZSU+SiLxJJyH0AVaLVIEKP+mb8M1bKNarIKsyxh+CWe4L2KxdYdsaaBc8
+mPOfd0PUypUCLdOr0OpyC3VhUQLHsokdAbyi/F7uPBlW14R+J2sXDCQs4JQW1EQ
nsbptqJ4r/JmoRXKCoilHAICCgHX39l0DkI8w0V6w2URMo2oHeESLwyxkCixQUQH
hqRZrKu+4zhQKsD86z034lG98VDQN8L4aj/xizK+ad9mxFgzR7Xk3uSbrYOmFxyA
48ArKPlaOvsaDLp2SEf320sF9ts8LSu+IXOpX0ctmqNE3MZPB3NQxqE3XosrmNS1
PFMxO4Zptk5BfQX1RSeTZwqCzZ1JWp6893SJrac9u+B3a1RDvji+ZYbeaCPh51Y6
th6S2F9Sa0T5ZpMrcPXzzgb34yAJ8DXgN+Y517qhxOV4S94v3lCwUl/wG12W4Y5s
Vvz2SHKls2Xg3XO3FkE4n5EEr+W5p7YgIj3nPYcKHa2PgWLI/FxAGRCth95BVMVn
lmlkCA0cTYFLOyVlj+bMEFMwAjW0w9ofm1fKIePYJHL9nTNXeFVpIEc0Wvd4bNyR
k2K26nsY6hjxSPSUtINPET5XYU5h97pfCu8iGdtNT9cA/hK3cMrrwr42iXX5bAZ6
y4a7yvhCUrEgxcFAhAbRcrU4d1nPc9bqREhmiz1YXSgWYM3a6MI0Fkt9bfm+Zy0y
MvAroUfuD7LTbwjd3jsjczyFnNf3p2btDBHrDCDZzHRClCafzfn2tXSmNXFUUv1g
IkKCWSYv4ClW51oykcfPyUN31MTDDyYVKnu8AC+Wq9MNqm6ZYaXY1xZ7BgpvSr4V
UQvnaj4jwOyhwX11SbwZSlnQtgQVVU9AWQwnJdYUsTZ0uYHqyRH2gUl00nGoj/8T
igeXqwxUhfFH0yH61uwcKWq/atPNU6eMnk2KVBIhWJ+LYllJWzL6k+FkoLZq3KMM
AkBexGfgqqNjv98UnM+jdrvB3zK/Xj2VHBzEoW0PXw/5ucBSmJvRawsDFQPRwDLd
JocjdkLzE67yNuJlhwKnGszI3KGba+1QETQ+PWesgP/3nvuEBj9vcWoZS4wA/ayq
jsAN8/ZAQMfDWt754Wc7lRCWAhqiy1HDQsuQ/hlM2X9tq9+fjS8CaM9r7Ojv8gG1
FOH2o9iIKUnjwKu8UE+WEsiRJKVOEMjCfQYPHD+4f8sQI2wRrBGTUt6RGefuAe59
bfA3NHAMhhguuSCIAqC/eh0j0v2reFGi0Zm9gkgskw0DejxoOh8osJgHWisfbJFr
ZS6Dd2c8TcJinGnDlxhVd0bYfWOYzYFMrO/wWbuHZFUovjQAWrmjh/rqECSK0LRg
cpSnE3xkQOzWkEOxdi7jbdQzqsYgT5wJnD46Wg2gftPKqscrQvYwLLOFizZZzn3Z
TDr7oIO5bl+3TbCeMpO7e3IsHXehIwOdx8YqMTHuaQ0JxKDLDF+2Q0BM0/xwvarI
w/NMWMF8nLPB2DHcC6ZeVmzvHreHejn/OtxfxXBCdUupM6zYt0SPwmQ62Cv9lqAO
asFp4jMkErLcQuxXSYlz1yiCCH9VOlyo/q/5CN4sSSUGBWHqSmUB+d+u2tFOOrwK
TNSCg7aLYd16FSSXaDKMt4oNGTAnJDHCU9BcXyA+S6BLKtGERjqgfkG5TPmac3Mr
1uRrQaD6X9HL65hf4Wg8N9RsQnWLBFBbeto9tfdbRc16edipxyy0CNLigvZBEle0
Dcjnxb/UwA0KCAYrbUjv8WXU+wYHUBZtuVzBjL1GKqaRQr2AcPD+H2VSvE5dwDEk
UQmUs0lBH13XEnQpMUhwJjzSyQmDCL7sYWpdCpz2gYyt/5yHWLrYG3jF9nz/kjXc
BLArCwz4dyt3XbHVtKFrqN8j7Ui3Bv9fDuyt+RBTMeafxcnXrMQr9jc0xHBpJPDc
0BDuk2M9IKQ+Dww4OOKbQYU6iyRxWfLRdjJ9RVv51QCP++L9Nw/JOuxTcLbrt3Hk
j6HD50sChcv3aH0w9q0J5BdEUN/xo9/xBP436miUO9Vl9x0+z1qFF+Xhk2CLyHBp
TpS+8sHmBsla4uUxmuvzSnpA9ONr8eHEhr4flnu/69xo+ZWq1CbteMnCXH5yf7au
Xhogs19GQvAMa0kMDwtrU0teDqgviu8mlaR5HhXpOP3WiMAvJWnrRwaqV3h7kaiG
E8Z3xx7+R9dSraDluJS7dq/dD5jpOFigq1XckYpVNaSKMRGKjM+RGXhZyU7uRyEf
EOZljEtlcxILsERofvGyNBBslZL6AtRvXjzyEcl+jVDCkvu/geOiTI2pS8t0TeDH
qfwOMDJbSOp6ntNr3bcXN5IX0s9nwOvw8uxhrgsomHnpCpjgH6RDRz31RI/FmW/u
STF5G/Te5eXUNnacxEPjlSU9bqdE2J5YkI3PiG+y2tjM7ZALFLO0R2BCENq1D0Od
A7p54Q8PQmcMsrsBrT7uuuOtv4uAaFHPlsy161eO1cbQ2i+nE5mR1bLDhODBrLj7
bYwXXrlE5KXAfJgtDXzdnSMXG/6KxWGzJVAQaZovWiknIxQRaWrqjz4NFDsNpA9a
8ZlUMlnwjmtH/ghFln+bAHiBU+9PF+k5bsCiOS/IHdudasDTULgUlYs8i9evBzcL
s2ad+w728V9P+mBVZ2AFfEmgO1rF0U1SUuEfGUMyzBWGo8CvkHHrixc/OrjFEqAt
UzmhFnSRKEaBZ54nBUR+Ul2igqcyr69BT1VxKdKER/W75PmXRxF3SHpzNAnz/pg2
yqJUZ7sZ0pq6l+LYP8EiZi/WUCyMEc9hpRzuO+x26jK26rTaByoTlWywoWXKffhY
xP2y8DnwWrVIIra2G+ms95GxonHPIZfwTn+KupWZVesslG5nvVn0ThKH6lOMnMUn
Ir1JD/CL2bUJ+VUeHd1+5/LSs57XF7vA7M8AHvo+HRRVqoQ85qBxjyUgqUV2Vtcz
C81ZmtL1TT/hNjOyE+hycgSd+mpymf3X5vhbY+fWz07njn7NaxUdy0PyqRepSY2A
Qx+IGZkudF+D0DHrkumCMaYaDZRgRHApfyHWo8FsE69RJWanPgOyEy/NL5YAsHJ+
5IqeCe6Ds7rqNKB7Ioxph2HzRHY6uibklfsClH8q140QwmXsdm1NnAc76CCY6hOM
p6ErHhDbPNLPbAH7u3Cm2dx2yRKwB7dL3HnlD5PfqJwCWsuzz1FvALA1KhvWGzl8
r67WvgVPXGXPtC8f3NDRb0b1l0CjU6LopXQzBODE0nRatIABKrobF02L2TucxV5Y
hK3vnxnu9c/FM0zfFHBr/hKqy4Ao/BEPL58NFX3u8CIFAnKnKswstA2y9PXMvyYb
TDq/zKwqgiGalqcfYgr7+Q9OfZAfdYYCQH0mTwBjvxOHKBH2ZUiLkCG9B2wpi4Yt
hzQGxphZYfAkarkBAwqp0ScUNC5I++rE1HbWCDTMR8vuXM/e1B+XNhM+eN/lcev3
cLyREQ8IBPHgb/uikLCVsxqdRST3oSY8TZENiKwEtCU//kUha63mB37ermWQyn2G
75u7gpi6Osp1U6H1GCxZ/OwSDZwyhAFGwnUlCze/0Lyagih6QHzZx1fG7XK+xEi3
GYp+emU0OCgiHi9/W4k1WW/c/+qzVBAMmNAloRvMGrzokRrv6GiAJn/Ufj95y/2G
R94dAYAPr63LkedtUr6oKpfWI1RBtlfvSopfCIySe7XC8NqUgazOEv2ptmbOBXw7
bxC+TTB7oHDJ8UTd1rY0JhzFRyw5bLKPoBiTiL51J4+DFB2nFT7cOGKPl0c6o6/h
T8Gc1pS2btlHEnUaoyHGY5deYBcsTi+MHj9JbYac5ekKluzRGhaGYBGLA4sPjIPz
hFkoxnu+89D7n1ta3Jw7XPlb8PPk4G2nRI9HZxGJW3v2umU1R9laRTBNcS5k+XA9
GJBATYgs/rPBoLU8D7qOKWjwazOB+HWY9Nzn7uKp2TAHvkGPmO3/JY95QI9gxODM
dxnlcAk6iDYo9igJZEYQFtNmBCYgN/E6mJA6Jz8Q/dX/+CDv3+9BNAuF4DSUmRae
5a1F24DZvnt9GjnatI87hPUlHrOBPJh2X6G5+zSYBUi0pdDuJdKVpd8MRol48AkG
QIG0rcQKO+ELo2u0cOXEwx0dJpSjLWvPE0h64DEICxj+Ay6csm2Navzk5THJToZz
7Q8nI/aHsbn6z6G/q64deEHWO9YKh9X0u+w4C1eOk3b87F2uKmmTZUO+TF2KE3qI
ZjxBLuOdOn2G3m6bTIknDDHyxMNz8ua/zJWtzYTqQQrnvHvtbRlnZHpwi7Wy4hQP
5uXLYU2I7uXGYyf0EASnuzdMEtE44ILTDhF2eYOUn7BH+nTRml0/8pw88FEnjW50
6EdVhfhhxFSK3atfsLhE6wCG6FuECSrhffK1rBQpipEslP9hTNLQNKt8NU7s5dgF
YgreQBwfM/TzFiXU/3L/eMNi31AH5suhBNbSm/QJ0148Bgj+9ewIQ9ZhCOPdHs33
aVdvi4/tbx2uEeOd9oOCFj6TpgaYSxLmFgOKpmGJ2sC4qHMfNgNBIqHoyZitlOpi
1fKkqZZ4vBhcSCjQDcJ8c8gcSN9BUVdH5ZGtKx9YZxS6ZdCaFzmyPgXraOBZyx/R
LCpTgZlLWcEgEn0iD7i2Y2Cc586imidspTYkzjxMmlSDb+yyyWxEy4ydwQVCvGZd
TAEF5mRGd6Nx9WB/hV3025Sp13W5m4lwziTsgGrLdjViu44NlDCbN/TxEPXBzKpx
OFV0vveDITJrIRzOdCD8GSvEnLlaf7+uerM0gvxeUIs6ls2rbwVhplGJxBDEJbHs
Ei7iVAk6vn3lkuF/aWB2+qY8+i7kK9/QxmLCwRjggtGIjIupvtsWFb0HYcvnnWwT
3LX9RTydOhA4S1tpZP34Dk6nDTIffsdLer+p2Mmhotir/31loSEmtKqdMMwXjXxY
Aa08KJ0wYexGeAX4TjmFFUuUEIj4MBmqSNlDLdyHx5XIAwjG9JXJgC5gw/Z4sR4m
cvvi0KPKVvSIsVvxDmQXtiyzBLP7LathRVgDVJ8h3pyV5y2Uy9ZriVN5SXdn2Su1
N56wIfup5RvP8cMGuaCoHxCpm2jcljJqJK7FENZOBusJzs6fsbxBFYLNC7X5VmF2
t+efYFGafQnAUxLSEqTzs6hOKq75ayox6yQHWyODlS1MhL+gmCnEAIiY58tNxZUR
u9IU+qLUdz0a5sG5Mdfp5xA7nb9uMrFJWaRqytSz7sL6/NRJDVLILFbNbWg7nrRw
9gCOzqy8trapvR2evpSaS0laGfNofDsbLrJUS6aCKSNFepOFBrK1HLhOIp1iiPjx
kfd9v8lfqafCBIxJxXNNwHX849MHi+jJwmQxKyOR2ToWHQgObhMJB66R2oUREw5c
690Hhlp39Bvn30V0p6FRrFUS62PyCNuej5HzRbCkaU+ADAym1/uLZEZOGAixT12Y
JjjnMKRXpa+uAp9wF+fpLImrU1vVk9scTSULnQIly0np0RgsmTUefjEXmm/DzeVd
X/tdHhZaDxnDsawj2aX64VWm1NW7fr0vx9UkFt9OVfrxukJe/YkICm5M+X/PDe+q
3niW37PI5VgMeBjkn4dZjTus7+MpLQwlV4Xi+yTPJV9glt3MOH4+T7/5zoYpcMPI
5KdGwzTcHWILz02NmOXN8oIPVHh8Gr0kXVqKwAxOM/1LJAfftmv4G/WOGCpZIgwZ
5hwrSAnOvDvjaJFw+JIKd9urjhKVgAeRpJjqX6sX4WzA7wL44Ckiw5F17dAnL24D
wGNiAAp6sRME/DHn/JDjyS0plOlfa5UlNTwMsqEy4sZDAHi4oZrKl7rwIpYkt33U
tkjL4G9sx6g4wTH5YtrCtp+v9cMY4Ap+uz3NJLxCfjHZSjXMM62jXrslagS/Rx/s
gI8SzI0qK9BbnprTI4jqkDqwFVmDlK3mb4QNvUWvlvAtC3yFl1TbKkwHrQNcLtCm
uVNPy3til+4hsnOjo2xXXkgdJcZ6spRU+ncBY590JImZMBEIVD1oauK4nwBe9pg8
YR6xRPpZo3n6vLBHoLfsjgbyW8dkiXYHCpVULF56OUTclwpwy3omUlGPKkNPho0c
ZZkY+uKBduT1R7ecxsBbTLZZr7zeSYzlyN42tCmFi7rmyHWe4RZE5oxGCrbpgzZK
ItkBfEzGUjMn8PIM+On6IzeLO8JKYhFbMezM55Hcwpffzd+eg5UXSXueOmmvq7kX
bB7pTVhV56/ZVDR/rBpWS33PCTl3zC3Om+Haj8hI2Gn35CZnIqn3WHs/L45FKtd8
pmRYKvtFf3p3TwKdqrw/r+D2NLbwWNBDfqpjjtARD3FVHD9N319owxJNtCHr2Tzs
9e1MH2XnQRmbSLfYC28UPrUuOxXv+hJezUTyhOvPkegLhBw71sEnjSXlPxOaRaBA
rFxkZim0ZnduI8H0HHXCSTYEbHSGWtrzx8tjS5oMA5pQCmJhhyKYke0hn//+kR6u
TDwK47u6rmvSU8myQIGtZxclZ8ng/pnr0p3loK4zO1oMeeygzFtbn/XYqHaXj6eV
5Fb6P5DsUrxS6DtEEA3vkUw01S5ctArIq9jiJM1/5lgTvUtHvStGluDH82raVqUz
L8a45WZ2nCbKuVsKuGkjCN3MmAX5g9dkAE3536UxRQBaygHoaw5KbVC2FUkyowKw
0KdS5aXclUOwzTZ9G5foWXVxqHchUzc2ohBbTsUcIvSF8eF6hXsbet05UYGBrNHM
339mPAh81UN3VBrHsgtf6rZym/GOaI6/sJP1X6SYvlRvSeyCtXlSFLY3qBvHkO3i
YDXFnsCqsx23+LGAR++mrsZsvJUp1Sm95zAgN9j9m6ZFb0C11xPQCEueVGCiB5f/
1AFYhk1i1swetBFWjbslmgfFy+hQMDq6KhmD0Ku/eMHbzU1rRQPYP/UF07ern34M
OXhKOw++A/5R63Y2ibvk/gE1S9aUQvgtdqjBZdBr520gvtWog+ed1tnUmvfCuX84
B6RRL7m6/qVAOsou5jZIJ6G0eABNtbgETnI36uV4JiHBNCvj57STAo32b3rDksq3
mekfoRDxFFc8DmcLPqejhoLBqqDouGHiyR8qObQmgZdZ3Z+TwbFG925ssVfbO2Lb
zTApktZ1k4JsJghavwJXoLN4neOmnGXd7PbHC06r6xfOsTb0roPjxGH+2SFpdOFo
L0ZJoiHhPWubmYckvbjhVTufvigHrFMoOKyXI2VSEzfUqXAtT1RYqnzFMMHOx6m3
AHGL21AevtnsApgdGAGouBkP0+efaZ7M1fuHfVJe1ldV6VAHamdTKMz6fj9IVI4n
z9vLs+sAoP+h+HQIiNdLZoqDwALZj3CBN7PsI6fw2AxIZiHBWr/o6mRLZZNSXrb8
0jFc9T5CGrXtmvIhFzhEmJ8Zf2x8JxM9vcByk3Wl5HO0Nlq8dugb+2gfdM/KJ+6P
a0ze5OZBzXhZZBDbJsuB1p9Ujn7skQWWJvGoWb0gkt4v1/6qg5LcXNBOTZJrMGei
cD9TnWTiI1SnCD5EK4fkXvLoXNzBFpn5RLP/d28JgANV3l4QNjL+i3QHdDFWwnVs
jNSMRfU77dsH3xA3fbugVErCszVg+s2pyfkvaa5yHErnsf2w2SXhckhaRKapwYOv
6RmamIpdpAwRaz99qyhVNNA0pVOJmFhSqC2r3TfDvAW7jtNuxNwCTsTLEuf4FIA2
iXl8zTDoTwb5u+DnamDoqtE8JT1iOZjbljYLySbUPFRkEmqoNitFetdFR4eUVKa9
cK30eqXIQh2mcWgg20C3j8lDv2RREEtRSXb8PMjXcjcqMnOGSpY6kegr88qd4l0+
jkbAbQ+dzizfG/MJYG59TEvdPeFDW9LmpamTcLHmmSZWvak+lK7evz1ehtiW3HUl
R1ZUtIZ7vmLZ4BOuQ2GdC7gcWixLdOj4iIjIFA8rYIc3NxsjbOeztw+gWp7YdiB6
V0akfqxKkdFYPzxpDqa7c84pGheXZg3M/A8rsMnPinNIUQUSphk4y2Q5NFJ4v7DQ
PXO5Dj/ZHQ7/czE/wtV+WNNlnZr7Nzm2rHxF0W5lbhfH55cYYKrGJbxgzK8USEIE
Wsrxs2OgSRInxBTbmQaTfYnLuxTQ/ZuZ9UdKR+8+XhQwbfUEYFY4zJqbJD8qgLxL
3HOrZmexT7Ps1INyp0EA3tuG2WdYcMc8Dpl+nZNRdifaBm2fybYExS7xv+vHHhSc
AbvM2CLoiRZVQk1dA3JlUP2OtI3g//o9ysIjjynwUdSGB/MPNKZbKcryvlUXv98z
nR9dBbXXU/nKg5DICDu8Wf71NOVzA5tBLLGF9iUJcr11TOyDVaISsk4XACneV0+E
r6j/hmCLCTv22AraD9OvYMczRUWZo0WK2AXD8ytC5sUqv6osM2kAlHBYEqL3qQQF
eb++Qo09LUCwBf98FEfmWWHrQUQQR74+goD71FfYfavVThYWNjAo9alXGzFQoFox
QvuwiYj4UgJwrMugEFdn0dhM+y49jHeZZP7ApENA864Nh/WKasVOm/TsV682Qnzg
tM8dxLcFj9VCYrByme6VSGjR76xBS3Ac5Kzqgmgo4dQaS2xUvPmYmmSmrq0Hfyg+
Ze3XnSZoW2m3Sn7RsUquGBVvNhvSULznIVIIkXcUFE5VqY/TE2I3eeoGpaPKJYOB
uCd65KkJ1ejS+Fzfdez6Px+WXp0OZXFLqwQmNWQSLgDyCmLFmCcvTimh0KdCAkS7
jB2Rz+F4nZgIN+Jy3WgQg45MN4buSHsgi4b90UCWcHA4eoqOvEPLknknDBPrXOA5
nGBI4Ikz794GSzRx71GyV1KuC4F3Erf2ex6W1TTRYSyVU3WQ53ZX3gU95f102RH2
gPU9z97WpjwaiGBj3VC711voOWTF1l5jdt74I2z7u0ex+NkIS7/JvMKZMafrxbFC
jKTRPytb5JmQlJP8j5HRhSaZJOBuPIvWauaeoSxZuDf0GJEZkefYeAZ09NWhq0Bf
g+uOZvgxV5TunLBIuhIbVMTh+ZyNOv6ZYrtsyu0wuqQ6zvF302DUQbNR4NOKOqe4
fp3BQu+DGV8h+yLbo79NtR53XK19RWFIecHCJQjiyZ/Ng6TNXovTnGhMvk/dXJSz
i7Qom1zm1TgT2+RKJMM/pDMxTNkLSR8ZrXKNAW1rTpyVZl7s+SLp5NkbRQ8T2D3p
HpYJV0XBfCCLutAStxH4Rg136FF/8SKnGdp5upblir7Meo1tBxzMqUdLAvrXaJ8S
4Cmn64lEKrvZaWQnKLHtqTOX136FC2o289NyghvYq/Yg+he3YMzj7s8ZH/ES2DlO
ycf5ILbUuiVycd7FSD5K7hcBUO5h3onxU5TNO3Wxby9y8DG4Z9ftqCDd+Hv+I8TT
DuqeJv4lRhlBhJWuSouN4HugtHUa3hbci07844M8oq2fsrwmAtjvDKHm6WhamkVf
MXo+ateJLzKr2RJ1iSF9cM6XD/tkknjQq5uTr1S0YUshCuglCsXuWDKfBt7cWp4R
on62s+rfLAfMWxQDKXomjQiF7bB8UtIrpMP/W5oO/wB90NryL/4KwAF9kpyFPRp0
3oEBGs9jOKFeJQIPkZguJEvu6QKXaE6kNeOTjCaTFHsbR+VE44r+OHs1ChgIBgTq
qi22kqIfcI6SMOuH+8Zm36136k+ji1g29uh5wbqy/LgoV/lCazsPOF+lWXLttLL+
NpfD8Otc/v1N95SuEdmdgTAucNjzEpFs0UIPV2+GXJCHW5+cLki/DfpnAJ9ddeTW
BgJFmTFocdgrkM8FGodl5zQbtFvdVOtqiWYc2KMfX8lFN9/kT+zymMXxqvIleIe9
IrxT2ibH0aBdRKj4yyiIOyl8N8feWsDTEOotilMxp4Sld3qUGwwpfSVQ3J4rdDgx
wKpc7U1btv4bCMWw+PwhWeAIaNs9IPpHZNCAuOqOqi0cwJLMstt37QH8bCufu6uM
0EayyUhNIOs6jhRMazaajjc98qcEt/dWgHaU1ujEBIyfjoDCU/+AG3Cq7wcxkopQ
+Hp2WNII8lViByh6Q49QaBHfuMDrm0lOB0NPu7miD31aadxP9QIUe8vsE2HtD1Xe
X5anUBDEfOM2SDKuzFQj8MagIIwzj6j+2b1DSdVzwnpcdnVwADkDUBL6wMkLUWzu
1/rLOCK/9llK8ivnR/VtFh6SV3YdaksTjA5BSiQsRTBjA7GuzHBkDLgMq/V8WFA5
Oc7ILYijnS65N7UdPfixx10xL1z5wEPwm5iBzjMGymCt62ZjdPkjlWtBJyCG2uYW
1uAh9oq3wBBPAGi1SgwcjRrsJUj/1JYa+hTbDYvFgDZQX3DIgY6MgyiU47/QLOsD
RLSha8+tkx0WKbkyFnLsvBDA3OM4pFhcfYYEZf7/2zJrHQBSAC7fe+WUvMfRwMmU
7auwqjyqiEHus56WmP8Anp+ww37h021P5/4M20FBj5Z2DbFeuU9y9lTgwsBcSkMC
ifmd2EQchXQ/5bbnxKtTIF8E3Tnt3eiplTQ+o4CJXzy4Tt75oNkgCJAR6WPw45Nx
aI/mgNi/KgtoV1yQW/MjMqfNxmlvaffRUuaRX9ibJujaa5D677lG2/l+DpsWs3Gy
kOe6KN5aPVSFeR3MdEgAbq/PHbe7MVmZ8EUVLURsb4ebcTD7e20BxJa2a/vTIHG8
Cp87Fa7psCRMeK3aiE5AMX5lg2hmrzW84WL628vPr+bROlToyqeHyuOzg1OYKf+d
8wuxZBzsScjnN6xylU+Evg001q2pvqOGW4cqMJ/6DONRqKG2zSr6HUJFjRo+i/tq
l3iDQLRLTNNNCd43wEhYlNNVIBw/j2RfBZz5q0AB5lt5V2lOm6J69AjT0s5xMw3k
sWdnBNClhGNdvYYXXg2UNZ5aKWIzaa2oZNYCB7y5aXqfSiv5hspH8/KATg3Tey3N
U6i/OPdEjKVRHYZtUOjhPdkY9u+8AjiMzH48vMh/5+iXm4Nfi+xrt/jmzSQ+WK77
RZLPgagBZROnY6ivqFNImPfLzcNmiXayU3OJ3shTKY65Am21no5a/zQ6maXaY146
DYEAzqw3EYes/dx7C5NGk6VYfTezuxzaXFZOlluvjwBWyeWgaIodBeWybq/kAH2b
5nmYPnrRnXbGhoAmGnrJiagRQ2lMGUN9A1qLAHj0HEPXO37KM+Q0C5FAUTqDJRHg
YA1NuRgJb868XillU4fufN9gUmrJgdJvctkRzAO6vH8CGgQ9T7IVl6K4fuh0whaj
M5Mb6DdCH3gej7zL5VDUcy3QfB9JQTH3+O1X+p0BhWHW/t6tmVM11E3Lz96vV1sZ
fo7sv55QhbR8Ts5utXp59kLm1EsIlVzZqELntFDFwJsClQfO/q1JC9u0j+P2MqU8
Uc3Xd/zcfF9LG354iG7RuQ9Ab0ZTV2sFggYjmiIUe7EQRSaluy5mofoRclJWJ5Aj
qRGEsYiVxGbyjNSsJYUriUXHO6/MJScLe7xHgrunh9uvq0xAIgHHEpldJBojH2rk
sMq7ot9bDjF5x6q2HAlHkldtTDmvJ2Sp0VSpoZpRucAUYFplj6wWJbuQDngdDV3G
/eE/wXGIszhK35rNUmOSxOtbC4pZNQZAuUswjFf/XcTAch0kWT3AixRRkPKC3hB0
yqtoPHLOnunkuOrwTdGxS294vsnhe3bmVST9FB7on2Fgo3BYpjQt1e6qTXzvbwCV
WeukPLwjNMV118VBnsMKuBY252TgbDLcbTpuiFVavOnmuwpvlaa/k8yEv7JzkL4Z
WhB00F9c1Me6GHtdBujC2aIJCbDkqFX0r8VazRviA7p0mbGNKxwML7mcXfLmBxt+
DFZZL8NukojYOyikb8CxLvdvbcgQDC6M5gbGVcEcXWqQBTOXt1DYVfu6g/88nITD
C5quS/WdIv8BkrgRemtLJ7toSJchMcjAUftT+2uzovi90zG42EYPt83g+C0OBJrn
ILpl0wa1kgU74N7sFKeX98LoYEwfpmBz6+u8H32vBhQLsdZkKsUu1vQjQg8oXgxl
eGZWMJR1C+RPtk55dWbgi5vG+o9bSpZFF78yjZ1towl/DpGUvclIWrNaV3XdMDNk
D2c7DjmBCQCKRoSgGBZ1u6HBOOeuLxZFpPBwxN1EKrHGJm0vpNubINh6f/7N5Hz+
nyefPpuFfBx0ouW+i82GHYssIYb+2CMImO02YzlaSfwKKW75Le4wditkmh2HSv5O
Hd7gH9EyvEL0flzSNAbTBoRreJbP7KNCS4OpxdnEZsZ2kmpkn8wGm+Frg6xIrfZ7
SuQB4t26N65NL2kmMVTbuX3dFH3UT7N03COniK3CDeGucwIvcnMcOm29G4tWjAov
LV1niTxsI8W/mRPvkYR/3CRXF7USRWGCIdikOPk6o/5fvPcMys7w6/qbgOOYZDBY
vGxII+YrHsGZeVmHpacudS9dIBZA2epHTxxE7naQILZ34ccEqFd17vIadHWsgQca
6YuYkvhkC4GVkDfR9dju3ta85Gon4TfhLWek+gbtoENgKTKr+gid+rFXddc8fPXk
FzE8/15NeU1bqqD83hFtgliYG7Qzn6Sf9jkj5aVqw4kPI8+zqfIce3xHYqigmv6Z
1w52NMmzNcF/CUsmWkTiAsu3NRxtPxIaDbZyY//YXAM3s4XxhYsOfvgpu0e61Kgs
kKIKwcXwfSSIhDOoZMJHgTmZofR5y4H/8uuAYO14ULm9F9f/ueR2KgqYNsnQJQcg
fiA5wmSMbBxMbxgDYQ6KQMw8VTjNEOywSInpXbo5tj5oJH7wXOzMsn5Qcf7CVqXg
qBCGeAzt+eQD9jCsfgpTAB7mgQdX4osiL69SpkrilqZ7/IRh6ylD1EJsI7rCXb/k
mGjNbxTEABT3vOkpFI9TeTiz4Kwskhehr2RChWnuadeg6WvLbLdIC6jbWmJPFv7v
37FdBp/dZMPA1NfSEVPpMTKnDb0Bn/AFvikELF/LI9ZXYnGoe7hXwsiLn3nqjMpk
wGF8CLMg/Abzi7+6gVQ9ZInsI6h9uPbRMLzgmaXLtZ2Wni8Tjk5ONiPr3RzFtEDQ
I/y8UXgLuwty+S37XpUhnTlFbaoJo9/pzIa9t0MSrkOr5WaP9CQhKXnS/fxgTOKB
4yw7FDImqHuaG7NoCpgmLNCl7TJbooFftcSHBT4LP3227YR+H/PSCc2lByQPZd4N
o9FTn5Edgd4bom4K6uK7/c7QXd/EdGqo81Jye8D8j2zdLubpfRmLze4hblN1LqcG
Dpmso+ZlvrmvtUmsp13QKsOmuLrOXGPSMpERVY98+0tomTJPN/ZgWMSd/bnYfLkP
yPYUpOzcDm7A8K9Lw4jVzGUuenZDIrrWoIF2deoMMxjalGp6IFE+D1PMH2gDdY0i
KyNJE/8H8gwyzPlcFWplj7vogHtKzWKHEKPgptq9juruOIRq+EMCvTtSeq1UqyXu
jCwOoEtNu0ns0WQxJhCfC7cpNl5noOtC6GMfeaZ20EQRJf5Nw5ZPi4SnugzagB5T
Sn4HrChnres+69ando/Levi9S+8gHUHMyFwGTmZUbL998jTfUDHhWUE97dReRRSe
lOokfu6Gy9WxYyLammbxZCAsi0g7h6PASIie1rdB7Oqn9pHPwMcoufQX8N71Dk2B
X16KlHr5COa7uq/ibzJlj1o/ewPKlmHyPNLizTR5e+YY5IYqDFVZfo+9+wAqBb5j
dNHk3A4RzCZX3S+ElX7pNVutirTFiVvFacRJCBngIhNpCuGssSIE44845qkrIkdb
e//46EaBZ9eqy2f/50W3K+GQ/zlgri0yYoafVnDmdczAdVtfm81tQ8f/661ws0+j
os7ScUxE3ydPceEysOQKuZfYh/2VjRy7/p/v9vinW0QcTKflZgumvonIZXvq8UFD
m0dmRQMI5za22dKJxZwurfTYWOsUpRDs94TPRfV8EiLitGEe/kD6jQkpD+3vOC5P
eMdaGvTDOsMUP3URew8WjVoyZbUzp9br62s3a69uX/Nu8rCnGapixpeWz47RzW0U
K5N1TyEl8Y4GaM6MSR0/Br+5ecmxVp7FnL8lclVSWGUb9d+h/7dfit4EQU/GzN4M
vERUIxSWmOnnDkit8rYbo9KFYgl9bhTZ8dT9vl3/Ots1RXJAX4pQ8G9YupA5FExe
Aklaqz3ED6Rj2c4HEij7f7mVgc4Se/NIbdWDwYvrmt6WPA7fmpfWKgv0Oxv8ljX+
fQT4Ve93Y8k/06+hIdlb4JXz1p+ttMbZiK+0usmnfG8luJm+eG5L9PygEr7y+RWn
5wiI0+oTfpKBUSB+K3WwTO/dY6zKmNurMcETiZKwDqPwcvaE/jJtjIFUFpzf3DdC
QM56auE3YzvuyuiJZwi0x3X4h4tNGRs/CsYTHqluXoqrufitPmUtbZ+iVdMaP9In
cBtt4P/nmLbKdGocptrCCBhOAXax6nKeRxL2uPmhDyj+rnb7DEU/zf1KRifAgqyw
Zs4Y3iN6ZLILshAtMQH+FIZXiQatJ0i7tsgh93tFgbxRi1sIMQkVAe8OK7HFJ4U/
FcyAkIxdK9L5NM8rWaG3WNKCttdcdBmoCaKFtZxZ72CabcVAXVIzytaDtjrhBNyB
4bl0YWXWObrIKBtVsEcJhlq23JpWEX36LQSLoqT+93fUTUosf7xhAB8R9GSK4Vh2
sx8kHbEBSzpC1VrQMTyZ89Mb/U0uBd666E7uISjj2xgZmLIeTeqFlQE2rlcOEjKy
b6dsQFPgDizRXJSAcvOz72Noy8stAZw8ANVAan9dLcQW2pIfv2f1+vXTDqvPIqux
vTibIlctkjkJiBG7B36C3wO3zrDvfVfDZrNzjChhycstedR9Oom/pLDjtWfJjWlu
K0Qeu+9P62+MGjXWAd1aj24pn8pDMlFc6cWwD/swVwsqY6cDJ1Y7XhQIoMuRvzy7
o7Hmi3MJiu72oGS5a+TKt9OTDtwj7eUFOPU9ld297+xU0GE4HkgjXbpdcLUYr5pj
LTS4WUfP+riXNgkpr83w+oQIXQPoCik2avw+TajdIdHgSqCf6gH/vRDeTvid2AJk
hR+/XkYLLtEqWW5odCsMv+VKSFY1P9cTlfayK757xzrz12M6//rojEH3xpRhaoDU
a3IZK+awRA7ZfKPmZxvt996iALpmy0WZW6zSZY3CV2hMyTi3Hc0Gsl2IoYpTC0eI
JpGTILLfxbsVV3c7RCNyZiVX7Ijc3+IBXmcK/f1KRSMIVYtSna2pfQ4BMQ0GYjEE
mFbK2E/c1BZO7fdiGbVn0laM6KtzsskBF4V4fLpu4r9p60ZErG3a+NPPoslU7i3D
OPmBbMTWiyaXfbf0VEfPAKVbEPLTygY3Zz+m90OiOYntVxVPiKz1rACfch1llTr2
uEPl4wzaApFIUbiqKcvEcc4msyXIt3FYeMNqpP6cov12XeHJiDEAEfYjmBIyGhyd
fhWwrGS3w3atUJ1XaRUwzoyHNP0gCI99I1Xiu450yJfVkclJpyygBeHtJz4pTOAC
ScUeuwpbQWE8icgtu0A8o0fy9HsP54R2xmC3JCnS4e5oShBerLD7szOAOwRh4rMu
3vksBlslxDVufx+kLz519VN8lYdn639e7eknoMiOVnMSEDIkfhcvb8CTBr2nrg1Q
5cKz2k4ynL0T3KpQ4OOw/1uZRUeavWVcVFU0hKbJ8Y2pQnN0s2/a7skakWd8m3Cv
bEkgHt4l5GMFodC6HOe7URa5qv3YfigY6qundvJv30yBxuAd00mkL7Z760P8EqAi
XlufN9vqLPMMp9k6Aragm6K+vuKIurLBSYwukaqGzV7gmhuSOcP6Pla5gcph7M/n
N2yc+AjhwZ7bxJsAcLvrIcuBZSA8K54ZiNLqJhn16txImBlW4IZKZDLjJ+3YBcHA
mRzfQALwFjBZXUQRQkGN8Q1hyAqUBEG65Y56kLP6hDe9rbsw9vWuFOSi6lg4Wemu
miW5wfdE+5wI1ivAY0unNdAaFfBfHblG8rzdASftQ3vSisPqiAwsAiKHU16Wg5MK
aYJ68iNceI/5Ue3UYRd08kfO8CXPF15hDtSZBeIag1QZPVVNp67YIuSlmaTKh7ix
jL/80wN5tKvUpQzVAL6Cs+yFlS74PsSsgYDgxVxAPFjQQdslu2ivu9gkXe3Ug6F0
hZozctqErhjuzcscSMuZMYM/9TdHhn1uUISn46+2VU8+NsAnauIBMJuONOOg2NPa
gDiRVs71Mm5rokwtEdGZKIvSktmGIJaYlUbEHySgPy4h67dDdo5I1etg+TgkEDSR
5gjnKWamBfu+iXrX6Fgtjx0kjR3DkpbN2w6WmnbK81UxiTfAh1nO6ljpRa2gwqWR
zXRdRQS6LoYEQ9Hr/mXmER6e2UAatY5KBLEsHxpzV7lCLJwWCUy48w2hDrlNBHbC
9FfWe8rfi04ccg4wAHedCkQU8nDgQ4kVA7nSzaXaBaREweVq6swulT1O48b5W0Yu
nme6c8HOdE1xyednUQW5KqjHWVFuxsRj1jES3Xe14CUaIA4VPPzWCW09TXy1VN3i
jxqJtT57yqfoTZ1PP0dOXMpgoaQNVVNnyjiJiUx3NtOhyJAYV5yjAdi2CGw1IFXs
CWsp2xOlVLzXle+JJLtK0U/HBJQdL9al+7182DB/4y5y6QFQouIbeaXB7dk7Gj8T
LH/UUMkyGV0mdvHflLHhpPF96WlNSBoEY74AgDoLENUf84BvMuKwhsaO6S+booD8
1Apx6Rw20GS/3FA/uE9m+0mQnbSKin+Bp45GepshjECwTLN+cXB6WEGpPslkMiyw
Dn2UtY/kY9aswHeS8B+zvs0+pcJ3THXTevFXJsimUtUV8QFB2DTLhYAHP7emVd7Q
ZrGzV/I9EYl1mYm07NqedJwCjs8MW1uBASKo4Ms5Ij/jlnffAMBntFMFTbjuYX5+
2d3E82Cv92CUM3yJn7XS/eTq9DkQEfBSU8WhagjNkm50oTvOmbPUSbglAwcuaEdw
pceZXk9W6Db2fGRO893OZ/Qnm73ObxVMYdAR3VN5pruklY/YZk2WE7Anb1YNGhof
JretfTu9wj2l5Dmyc8vWwDfgAvsOiis0rOLBu6EFKB63k9p6co9zbbAs2/y2xIoc
CX2A6IORZ/GDlzEvqwHaFklVjPoyFXRBg/dn5rsbc4Mat7LIIWBcvcuo30PKRY5S
wx1JVMHkmlbXuRHgpRCchPlMz7tlqTljqoUtS2Sp3aupfkiV+klaEQ4AGeWOv0rB
bH7HXygjVQpp+DHS8CpR++UsZGLna146QYOtc9RpTM+7PeRr8eftjjOrQTprXTg1
cW50yunBW7crRhFfv0/nfGiIkR0ZQOf/hQRK30f/eenjIK4c4NTP+rH8bSE7rKin
YEs5YwCyy/OVmETDbiFOFu3z5GrNzrzn9QF44g8HXUtFrizodsftU+oAuxjARjr2
zM5qWOE8FiYiFFi7WZGnWqBr4azx9AfunbqwGgnKnPBP2KUZIBqSlm8TRSxxXXXb
yvxiKRMYAjuMKtV0uwJN7ss/uisMqD+Jmm37OqGF3otuR5LsH9i/wkwx2LqjIBJN
0R4d0UYbhqcAO5qajkXr2UslV9pxRabL4QnJrN0NT1FR/6Bz7NhhtNfimLJOxOEj
Cz7aojV39LIavCzJ+Ehblbe69lZYv8LiOJaJ1MtM+W9fnc/IcBQQSOlZ7b77+t43
KjY0CMguL6y1cXCiOs1hhoVTPYgZTKWi1nJqGm8txsD9XQhoxgDbUylX+nZwawCp
a/CtYbTuaft+vWf13TY82ScG0y6MelDz4EnOUyssJpqsbp5UWQKDEA88nGDkBCKU
OKWOyb8jmfqsMOi47GTy7ctUlosUSYnrqDpTve/9vy7xbd9R/sRRVU/iTw+OIm+j
Rb/QpmIIkbLbLDaC1zY528xv7bzvDJK+A0+t/4SjycHNAD6oBPjb9ijFsZ/R6WYx
fI2mu16JATfka9lIYME9fSytOf5amwbIyupo8BJu0K184bj8EcBkOldlvZJ1yaHS
Qkm3Qz9afG8+E+zkJU0UBSoJVAvDtoWlUDv5NsjmrtCZ6Fzh96ekzH/GZUTEhfqw
VlO3xauPvWrli5O6lh730zn2wVxqUST344G3JSoFv3SNj3j0UigcTiYwBHC/BaIB
fX2Ogr/qeq2UCoQrkcQdhekFHQOCosJlpWdd+aW+VVYJh1L4MAkanm8VWaIT/cZV
5s54kgMg+t1ZjlOkU6cqsmQgvPaRZ2UEQM0lUXe4RGgrzypyXmo2qWi7K5CLhka4
Z1nWhJDSCloao1tfJhf4QOjV1m9PCwbdOiZH6mY41XjMzbjbxHU5HtIvQYob9MrB
VPgoKJQKpld3ti/jaiiVtYQtDu7z0gNyuBQ1dY5LtT+Z5F+Y7X2Qideq9ndxpvHD
eLp0fryyBnA4139V2yq06xkb8sVfcc5rCTcD66PJF3CQFkCuw1lR7gRK7skXKd9q
iiBOfy25rh/pCTKCO5OBXU29NXDonghN++kTp/JNBRYF/NPCoeYuEt0iEzf/bvIF
fy6maIv/FKWZren3cPvHrfA+4IJRGZ2F8xQqYbfgGGYixwZ3YOMHbCBu65O+sNiS
qvBcPIoNDneX/W+rR3bTHcrgpsgR1UGwZQAapoOyBGyii5Ri2l7ne5SBeZzoEMPI
jq+sSAKQkZmsW/zaKNb6GJuc25vkGf4rxEG3haKtTQPtFM+3cgQ5H4f/Tor32qLJ
SWS7ni1Q5D2unjaIV+zz6guQszHoiUt0gAFrn0tn+xD2u9910/ZYtkTiA12GXeu+
LY2k+GVBTr7icM51mwdY5JYkpEKAsM3nWv5Wn4ZSrw5n1Zd0IuIVj0B6Q/USzDhO
bvrce/SFmuJYwHNXncXgPxdh3qX/gLX8EXW/uM61h5yqpqsmO0zlAjvoEIta1447
/zogN5pvgYYfeiN8UcZ/71jI4aCroZ+tVE4bZI/7SMqg9fWRatMJ7DYO9EjAoZ8E
/J0c20HRNek5/QojZ/2X5q0D4bXIC11UdfXZq4Xgk3x+mKj0rn7N9o+C7eaYxzp7
yBbVzO82t/V3/UFIOhhWI126jaYeDhRTKqBDe59pUEBEXCea7Y3bpZrt5y8K4n5D
g37l95JKehkYZxu2+KQ+SQwi/VwplNKZ99OEte5tvjxqWwLcht0DXGhI49CNGufB
hOCtEeeSZ0huHlUoDfpd0pPI0VX9UwiB+ZEe8ZiJGV7KAh8XDYzsz1n75a+QuYU+
RKcgzMBAe55YOqjMlQaRrpogvGVcqMmIT1JoMdHbOXQuTrJrCNYzIH6eN9WaTmfs
uQjq6OG86JWNEEzdpYWuXBVYI63fZe/3fhZG8qR2sduRHjglmc43vxaUCAxEVqWy
7uay1u1xqFjSDa2fz2cGFj//QUHg7ujB/F84shJPxE5YF9JMi1IHCtzPD3ajbjo+
S4motOSWCHex1ErK09DeCeg9KDiBr0sEPnaLHIG/QWyFuB/G6uEuyWf20SZBgMrx
NlbetFURmg4ilRfl6ONdpSKo1gqgPBJL5PeC7FFGnVqLjKwWYlIKdhzvd9Aqdll0
hHUE7rVrQluAgl0ubiccrdS6aaJf+LpNOHRy6hp761CE9s8z/k4MlteasMt0tgPu
0ihwiyS7bQqsLYKQeL50FzOle9dCIjMtywlgq3POoWZCp6Bxh4fGUZ1JGG3wNBbd
whrNVTlS3vPzXpYr+y8Go0LEFObhx0DaDSf06EpjglUeOnTchLmRJIygRWzxv03o
6hdrMuucEwK0YAstjWwipQxd7P9LSNDTuXK6BeYTr4+VZIgcIT6ltHA6QuWI+KDW
Ov9xJG0e2pyYj3EWQvmFavIpwhC2fnmTe+IShGOV9nb5Wh02xRzYSdCUmbk1WtiT
3ou+AcsxUjA0x8CNeBjcuyAxMhLZtGiVqA+gxRH6mC/LFmYR/J2T96Ix6/5VpnUN
lp9xDysNLngiaGHOr3qtbRRDlxRjHvHZy6QkWVASlh83nXAn9BXmU1tQDWZLcyn5
sRDZpoZP+C9QMpF/9ojX4wDI3hmLGkmq6LAQBpzSKM6JVdYq3qeYiy2kH+5pKu/m
k83i9vIU/JlMRLNvOM8Eh0OzdSPBaUHwPbvpJ0np7PuVwHhjqaFwEPftOirGhpsa
J6TjzM69CgRL5i80kHd4iznLNbsj0dmU6gK7vffO2pXVphyMj9aJjUtT6f12Hsiq
fXB/uUXYZqZfaFFYP3N52kt5r5mcEu9/yIMIAfwBGrLh7mKyA8EaPjuNVyhiRlNL
ktCMuhO3Kp6trwuMusL14Rqavh+099d2+MJg7JsFBHt19SBMpm4hd2W+P8nYReDm
ZFzerOGnhfQW29OwQwf7O+C/JyKDMnvMwG5Y3G6pbd6TwwT8fCuNod7chBaDwnJX
CvRBrCFlEQlYL+6cbhIt7f7rPLlzFGwMhy6OHS2Gt035p5Scu1oKVyxjUyZHVDMd
r23u9muCl0V9KjQ1WXHriA1FiCMx8ec/BAAyP2sZNI40hpIsqOFeR5RA6yFbG/HH
1VnHfAFqDzAu/dou2r7QUuYwI1UT4R86zr/L+EyheIJmSndFPmdLjKIIXxWjBl8C
vq51e5QO6qTmNRO2jnIJDv9uarXksUpWBgLaccxP/XNe5xmqghwmaZ8+y1B6TcTc
VZ/bY7IiAq+KYnBtcyL9YOakofhVE8yO+0zO1oLz8YDPRI0CwiopcBwqsfwQxaKA
ACYrleMGMC0cNkuhHXo8TZX8Y1bzKj6B/lLoGznG3yHpztE7LYL/WTd9ro/hSy3l
0BHraxn4HSiodQBZs2EknfJDNj8keSfkbMbaqh7E4daYBx/UjCemnbxwZwhQb8Nf
WkFHl1GCbnGewP7EaQXl/ydzr4vnEITdy6Ou8R45fA06XV79fniiMQFMhiA7CemM
ngRKCbE+I0Je2hw/k8/01erlQHbJgh4aSvNbeOQtRkLPCL6QmUonYRpvZmRqR3PR
ibjyXlDzqEeI3q2vqvlhR8YR6ZccliSrNt1OqCHj+Rm/hKpGV7yIClUfnsonPdkH
RzOaIqUzPiXwVO9Z+U+L7+xYxFaTsfvVjjdb//9F4LJXFCh37nYbFJEjGwyhWUmQ
mqM7qijDxwzQxZ++Pa2n1JOTWZYHbj+ahba9U4cpA4qsaMN8FklW2ygzDi/TeEKi
iMJMEoCp7MIxumHOB3K9/LD1qh9DfP52iqZvmspei8pyHGz3FC8TF+sBbCI2lBwv
i6PO3hreHpmvA3uEWEaw6ItPsqdgbZqbBlaZe4WpcqFTOOejIoj/ejRaujeW7Cv1
cDe98RTnEwA8eZAcgdVkFoRVXM6z0Bmo44U5FhRXFOk78/U056icMyEdUDRRNAbW
hOBa+tAbiVYN95TyQ2Ul7LdSzuQeDCOiEFt3oDi9WNJ/6Rig/0ftGHltNqYJ4qZH
+wyle+FuuEpB1b/zcmYIw7U0JgJk13te5NQ8RZhjEZ6oVZ6mjvSjGYG/xzSGQHU3
jL/F5d8cBou8H/qJtS/IsmdX5J7XHcVE9KMEdO0SuRG87FBsOA4tB4fRWw/j4FnI
+vEjs7QvYiuw3glEgvlyMXBaxn2DMznRyGxjBG1y1AJo9yyUqFWTuHlDPMwNI0iI
UwRqV3YTh7HQdBH8VIcSGD69PNsZqUplS/L1ni2YpaXYEDtc0xkjKs7mydbdB+WF
jWm2WJs6CQuJpAMlCmITciv81fIlx59djC6P2QMOqp1BDtNzmxbRGpnhlOZunPlE
Q+N8KNACJGLp/teHOiPaC0mbHgKaLo+DAorWbHNgNYCU4ZiBMIc+Xyth43o7S1IQ
xk+4sODOjxLOTVQ8iSlEkqzhRxbD2uZ2DRMOWyiXJDLK9y0eSN0xMxr10bjpverj
BXuyrhTaTf7JEshCW7FDipto6xKB9wgXNoZ/ajh868RdQ9lY2CBnG7hNhC5nQ/Qh
RHyzkHxcYi3SDnWmS4iHl/c7ajK22VA/QKvhXKqIc6IHR+iPk61b9ilrbvHZVaNX
RQihtV7CHSnupv/acrsHEJyQjUboxFAk0+++A7Gl/xOStYl2qiox69mRyVJzmpS5
xDv48cmMcgA7iaEK1v6x7bDfhHu2o4LMDGlxKgFRtOMjmboF+2wKrZ0rHF/XOwV4
l6Yj9VOMWv3W7pYMRRTgosexpmmNwIwqbgWEm1Rh4CtMvU7dd3+whQv1hH23i7xF
tTsxomJpGMcsEGYV0gVlP6LpPWuia8KQkqIorMgz0/Ebc2mc684I2ZRZfFt/QyXe
VI1lbHakKznWRhChoCZDky0L7wVZo0Cj09n6buTFgZMlHc9GjBYnqOqlNjEzC15c
YD6tVXr0KUnOUpUT/kvBPeT1TdHNkp2uqtpBJAbV/TX+Wg1GhzJKQJoOEkuytcek
8yvFHPXDPvDkBcNwevIzLdJQFm3gRCdHDc/beEF2a/Fv2RsYtGpMNS7qiFML2b5c
zqJTWICyQWZQsE3LIpnz7q6g0xa0ZJJ21eMFP/jVSr9PURU27HwRTn47TJ1i3HQQ
Q9CIBxFlYiC7a+Ll6cL51tIldGeQJh6bMKZHMZcgKi3lbgNXSsMb2AeuDwIuYAL8
7Ad4mQgjSiPSgKyyWoVef6Efo6xinbQFVZfXsZHtHJ7wP7moqyFuZK3C0tD9EqOS
LmIf2jHSZZEbuCztWkjFOG3ektlD5jkbPfcf2Vk1fZS1zk0wkOqGyxU7JGd82UhU
4stEcms3vPC2nnqauwiVD9ucgo0aKhC8SAVLl4K3ncdQAENG8990zcY5mFWQGxJY
n0rCH0inRRpiFHI/aysaUeRZ1hboUWD8RpbFAJfJi317jT1oG/c9TYjfBLylsWzw
K0HpmxFjyGmPsx4D/qwfJOl2msUMFp+AphhVcCQWJczT0MSqwHAd13COyeyXEJTK
Ot/b2kX158LnhMUh0t01cK17A3CdAZOWNB5JjCBYIIYLAeFh3trwLVJqZ2anZWhD
julrx8Q2rnGrIUkpaNcNpKG3CEYcHGKbq9fsE4WO4ucSYrmrMEmSqa/HgRtKjerJ
O9yBCnUKnS2ohVNQ7b+867cSS9hXOO1ImztZnajN6SXiBe8/qenpMoU0fyX9Xo2l
Nw2eT3ur+6woEWhEfoz7QNO1Dr5PRyddWfWBgZ9zt6fcPeDyrBedGRCdqP4M3EUa
57fUMB/ayrAc1ZHlgbVvwr0k7Hx7tkq/0Tpe+xYgveG0tEwS2Y8sKOrVG+RFHqVZ
DYlzIxbIEHsEdatBJVdfLQ/88k9qLe3gr1C54a81JALVQCzMRiL6DcERFbfPqjsW
e5cdwTTiQx0iMXzsRLlVi06/A1A0DzegrdG7LjsgeFQCJELYWzajkkMVdSyHyqda
YRDEup0iwTZ5YnftcSDCmVH8cassKw/7+jF2qWTzarQP3bqz02r8wkv5HGuzoMvM
fVyVXzGykgqf46rr5OudGL8QuL2u41/h4f/GOanA/BzZuS8mi0z1uzWio/8PotrV
ZImTEe4TL4GxvTElM7KFqQdfqwdtQnpRrpDoxOY8NJBWHNcezkssjCMzIGicTnpF
LzBkYkhv49pJ2XCNrwOBo1zFBXQfLrjWjkY7daQOVVCVi534aWyMMqtyIJhYGc89
0ZBx/yMh96S4IcnXSH7FlENxlam9YllAkAbxDmKDaVvd+5CeaEt2/qoIlVYZnrgg
RA7OJJJbCScRBzJ2sKA6rw3SdK55I91dWSfaWIGPkcdwzcdPkrM4F5iazIU0O49G
9dzIcbwL1+MDUlir9zJNA+g/9ivsdLAzubDeIcuYXF9sFOKEz28aMXawflqv357X
Fg+c908mNq5sn7qvZceTkianaO6g/D6eQB8OcoceBbxdH3aG2gVZsm3sjKB5Z2/g
nzb7jNvX8ajOBpOP49/vu7GU50Ri6XCB6vCkT2FhfMarxnrcOau91Vhc31Sd56Nb
+V842j0jAJclGWRCBkIUgUIOGoA86BarJKkAUBdJQeDaloq2axAvfIFVEZ+9eqs0
xWXLqnt8U6slghK4NWLBvBgtCOwd1Q9yEfCC9aTB7NPnrmZxZw+kOxMers0fycv2
eYwTWft2+g8WNm6XIBNWNoYM7fDPtHM58/JMF8/EyPSlq6AHNFLeHpfJVpyBgqex
EIrWBjcvgcuMTnKmHtxatNDuBO8oA8FIpvEoRAIqK6aqbkaDiu3W+IWFete/sgew
ia/5SOveif6nqivecnmmhZcLPAaMR3odIp09PXL0BSHTo0iQUZKHlyZhBtM4Ki2g
ObhNvqb9oyiYfkZsNhrIJOPvsoVKbbWU31K/dYz+dv4+klo4JptoGZ7g2TSe8CSj
LK+JcfsB/1nXePoCDC5E51xbxLaJddu5goijc+QsaiFLZAaPP+qyhJEOy0dYDxM6
oPiMERQs6K4Lu0Y2uhLUI4DVWvmrtRNo9Tsu8ytbSA3fIprqFxrf5Dgoy6NUtrKH
8A3LgamroaAO61MuACOA2YPPKnjEq4C3NCXb1r++d5NjykEwgzbT/SjeK5mcqZEM
W/DAePVld/h7bVcGL5QHiClcSNSo0zN4Nx1LHwHhKfumu9WIeBt8O6WprkQDLcHA
gzzap6cpJsMVCw0kmVHZERnreV3seeQL9pucPA8PHdzU6/vzB0f/UGlp+3A+1js9
NpqisJxSFdF5AISvYbxjted2aHI6c8kXIep+LabKUb0awymED26TDjANyQ1gxv50
aOnF49GqLkSnjfY/RY/W4mECnFONGrkXs7cVAXKiloB6yL/XjeslL6+Qm0R2Z9ta
LF76UrWJI5R4Gi+2xrraarPXoALZByMpQvD5nsM4AGxD9XePQa93hDXFJFE+gHE9
emAh8Acls+00v71Hi/Tq4SEAtOX/s59nEPKv5pv6lXCz7JHx3RcOjDhDa7Kjd053
y3lA0u7+7P2Ylxf8wl/piqx9T5+Po7TRoyDArBKpestqrC5w+djBJ070T9Ea67yW
i1ACCV9WtwT+TnwaWvPQ9FcUz3pWCON/iB4EOf0Nz5BPLD9pG39hM6qBKhsQYDnL
5Zn3Y+heW2GbRxuNWKnpj+s5a7AeRUmBJ5Yg+qSX/cQ0TXru6mzeatxaPkbehZt8
ORJ31KpYmKI1H2p4Nl83LnZONKVI7Cte77nkAraMNmOH+n56fVoPKH28X5aorois
W6Aw5QcPuHuXAdsYAAtYqG41mbW+l+FiZc0KpeK/us5hmCNwaLbB0+3rlWt/exyC
KfVWXWO3zGWzX5IDg19oGtBSFs22rm3dQPbkMIxAUNt9BlPeFC6xYW6wPnbjhaVe
6H+oQ7lsSpcPXRo5FmCp5VnHz4bZ4VeIj7MdyZVoSRJRLjZGTktHGGZmuuLe08on
ymZo1B3BLxoSN/RKM6Z8FB7vVFvFSHufwQcAnQYZMyDZNAOIQ5z1+fl73qHXTJ4p
637nkvh79HpDeurGQMF3rPXFip6cdNklKYRZn8fOM7ZA3cotTnR1f+uEl9Wyt9C+
5RSivImuFThDIOsB5UdanT0VthVcWGwcOsBinlxEwzpSfUpnhWFI1Nzvfejm7wRw
yiINrjUiYQrvYF7T6G+ar7O+hUgBefxzQSr4SxU4e/sT0xMrwWWrIx1PKqtKg96R
eRQqt8+Mn/fZ+2J9mLkBmILl94iNdU/+DSsddt69aD4OWROqhEaxH6ZJ7vgGwsC+
YU0GaxXuHxieDWLk8rC7/d73oxCbLd5ObAGvJ3tfgPyEGOzirHYBlyt1qW0QZDWc
YE1V8Ry2mVmGB8T7BoXoAHpIs0FiKpuDYv2pBmCkFd2HjDxnqNMyJ/mSiADswRAG
ZdZY0pjBUZC+7yHpmJMVb7hMMYNFh4OywyGXR/jq+kXsDOyVkf4IBjsJASkiZbBV
ps6Z7aACqAqhizzvyqCyevMc+8Br8o+HRmqd81W0XemVOGC32Zf5snBLwArN0DML
6ICBo8KfWKQYhtprC7/Vgcohbk6iY/TAYux9/K81USVekkQQp3gatmIVyF1tQAhy
6Ta2n0F0OHQzYosEehR0pRV5OkLxziMDa/kWiCnezqFnc0Y14PzR9BsMJYdkgmoR
bB04PHKsUUonB+s/99eWoomfAFjNwBl7eL66/8VaoEqM7QBsmrQiWv6HpyHKRU9Y
n29OoIxD+2QC88kV+ObN/GDHFDB0oRjchJfsz0Yxcl4QhIgnr5FCmzyBlwTX9XO/
F3lUuo0A0V+vtor0s7vuRaJ39zcOa78MjshYhG6y+3lgCpzr3caHQxkuUeiXy9Ue
bHHP5Z6Hy1KUjnlk8qFpSc36Y8ziByL8tmC4N40TMMM7DCm0thBIGs5rTeq97Fpf
SIda0wbbfnMafifsAK5A0gQT+YYk7poKkNCWQMAdLemE5/g4owwg4XjGdOuXCHZo
IuvWgURyf/M0GnlbUMlhgsglJpJKzMZjIzX1qkNBUjO+8mUW2DCBRu/nIRZYTGAb
cxpNSTyJu5LuejdcUwY1NJWYvsj52tVYlLl1pUPv5wMBufsRgeq2gKv5qQf/pIu4
zSh0OqJw3/fDU/xUaFDpDS0wqz2zXyMJD9qrKdsjvhav6laTu1Dua9OSEAKA/C27
PB+VYRwK7rVVO86rVWOTrdaK51twHXF1PyMTa3/iR5SalpNOpz9xrjuK35c6Jc5D
duj6MYRYyrZAUVKGhBGy0bHVnmxK7fUMDmqgfW5wqnzHvFGGMxvi6SanyukGYKJj
yvRBAfWZKg2Pu/ilLpTzNxgws0I7PeAVIDZdkY6G6JyOof6JumX4SPSwEUjnpJTv
OT7KF3DOkTibi287pL08UYKHVZyiRKa9qEBEZviqEPYVpORMVJN03icDHFw3DKo2
/UGpJ1b+L0kWTSfdme9bBDiq0iQ44LF+j6/n5TRjAwE4J5LzeyK4ytYuFU9y0Zr6
J9/KdZ83r7cm2WV5KVrIJh/rX93dHHdP3F0RsN4x3zmQwOWQqij1pSs4zD7STtRW
KvXRXbe7GwNlylbk0YEDfesbwLYlsh3PTeTOBxB41tqOZS4mC3vSSLc9cAuF4KVn
0u5P95rUoakWYW2AJHL+7BMWw4GTfY2usKM/1Y0f7kTdSFnCI2BogmSeEgpFE3GN
35vpFAtaOE5YqC1AeKyLXLSO/Y0nZ4zY5Mhq2WYRcgAL2MDOXM/vSwpw96hzhcHd
1acampAvC2rMlKZfN2MxetM/MsInljwU7Zq19o8+rsuognJt/hr5Jrkf1I7cMrGc
RU4wZEv88QfflChfNgBv3Jvzg7mHON7qnVyEy++I7X5udv38NlAUeoKPVAbqkmPE
j6RrTmoPadynxC40tv4QjsHenbfDuY93yT6FvVBX0fjTWyQ7yp59ZzKMoZIhYiHc
SlXiw4xY1MhDSmFMIM8SPVDcuw7Vpin0ICMp7gh+yf3J/lzAqaupSJB30zzYkyCY
wrP1oB1I4RNEzd4id3LfPzgX8doS7Ju0jM7IPSVJz7N5IOgJcr1cb8guTJVS8WF4
figdmrUQG5ebkDgER5uLkoTjLlmYL/Ukig/E2V87v2Sv5bndmcSs9iI53LY0n5fi
0nBKa0Zz8EZGREb9R610s6ZQOEquQZEb6EWz9Ml1KARoj3X1xfQVpczdmYYpOS7r
MKByaC8HuOLS2DE/taXFIu1O9IN3Cusgv80i0byzB/QrCSfM4LSEHUfTXit2KU8F
kupOaOqOAUuL3Ttsj0C3aYdC8ko3P1ZIEHFyO8XsOrfeCmSHl9+FVX0tjMARgvxD
Pz+QihambgGOmo6d0dpVfRExDvrspcIlLXhOntbl5u9VSBn6tMmaN8sN0W4xecP0
Jqj2DlXMb/iavFg6uieTZ/gqXxgatkZLngM4h3PldoXgseZ7SA1GUBQqJXN9b0CJ
NvSNjLx2iP9rjMsyUchoeG0e5pPAMly8MGlb/G0NvwCHvubHgp+F+p/Or5/q8Yfn
Ftam1FWvkxQRB1GBH35fFRTfmlG41KQvna2euGizdbLlze6lNiGlJSd6XF2GDsn6
drm+g2bOuvRB+4RI9yuFqJ+vXKKLF6xNwKXu6L+8Ke7jbTWynb9ynsyxW3HSmke4
PDV1a0PSp+QkAMErFbyHEI2ySQ6ULy24PRtajtzq1DHfXCDiWFPIXLSYZ9JquXa2
E8Ya0SW/NggRPwGbOdvyRaxdD3Nmf7sX8MsncudyktSEneiQwks+2q+Gwcor8Yq+
77uurPgdc5j/Sm1wG3hYVfppsVPI2VRXKYJv2gUCaG8wPjgedTkm2xRoxru8HGqy
gI8zT47hxtR7a0woXLoqrZkMuxa8tGwwWTid/RQaHlIRHjA92iU7oSRgHosXLNsj
Av90qQNI0/GkT6elpiUiF+1FB6YqiEG1U3EXuXX9YBkp28u6cbZh1KuEWVFFPhHN
K1PXfg0Ffye51mvXE++sFclh+tgPFQnQt4gL9ZzfO8YQxs+wqkriP63swg0p5B/p
XKRhOaW8nEFteAvAoTt8mHpZNQJIi1EGWZWOW0iE+k3yyXoKMjzUEclYlE4c7Wj6
oAbE3yuo5jAqBdm0bgZnBd8tkyFClVR87KGDj2RYwfG62Kulh+qHwwkHeLpWzMbS
S42jacGmhx6SVxCaiTe0Txd2voe5sUm7e3mGSHBs6tHflHol7EWm++0cgP42x4gc
gSCB0BE0QAsyd903NrBBDoIjqegGFZQep4jn1zgulJJMMYLEvUzZJNsO4maGPedj
5oavCQtH125i3GGrMV5UNsfrrOJle24zmUM0k2Mu8vSs0Kne9zKSkvTBTormlhoj
OodT0Ki2vmSpAark00mH6s5hZPhdPIXAiWDcACQnei80kHoT46QKy/BghbTdaYxI
V5ZrsccI5pHAZyrMn1OGaJ95AsxT5L9L0cow86+OzkHLWsvhP5ve1OoOB2khpljn
RgwPqv+M1HSsyE5LLQqSsGW3gq8OmOJMcup6EJh/DzpJ7YN/w33RTaEJWfCun0OR
OmlJOej6xVH8ioULEJN5jBhvF8k/+6w47KV45945fURxPGH4uhkcz3N9k5vijDJX
0Jzo836UHlYGY1x0pFkQ2H+jkJqsBFxaNqTHXsGblPZlyUXu24dXSWTUf64xbiHZ
30rKwq5v18wt/tFO547QnjlYBDyZwIR60w137kU9K0k9iKQdgFWjafOL3AQGbvNK
PkdXqA3eaFU0NEg7Na1sI67D6wy5GTNcoxgbopDDJj8yKKA4ISVmFahLBXOLS34F
1P6P8y/PuKUopxFo8nm56khxV517AD6eL18yKV6nwZrAQRHwt8vW6TxY9JBT9ENO
pGnRuW+4hvvW9Aazo1ORTqHmsJ9WMRG6ONhywh8A2Z3OEKw+bEC9o69YQxHqiDz0
az/N1sHw7jwaUDn8pKHK8jVRK7KnX5iVRGk7bfLo7tur/Rs42XYOw7spRj2OSE0W
egSsJS5m400R1IYy6mZ6uxBUC1wfDnldwoRNSvm/DBBTtWz9ZbXe4KrTjPe6nKHo
tIqejWyFUAZpiMidNrcQm9bOVbEEuhlCYKyx4936ziWKDC0Rp0kQLnrqDmEIbLzg
/3AO1jVDeHs7VO0tcrmQHSEfYTq5P0KT2umoYgSPin3sVQDYJessTbVyc6axnz40
n/hd1+UY5vcOpCWDeGrxSwQI6Yqrii5hc/1xVwDRxuiYOT2/W5i/BWzg5qI/Ns/s
6ZsGa/v/JSJlzoobuifxFjYIYnhaWRM1hZsvLy7AsWwpeI8vW0Fql+mv5k8FxYrC
Hg50KHUDbbEn2KEsR+wOkTZgUrJ5L3kY3/+0rYnqXR+Sv2jQPQoax7Hs6hZixvvu
dDVUxt+PyN8KE5Xm/lKtusEgCCZE6AaZ8hM3d3P/bPoRA+wjR9e1oMdkodFntPSU
pn7TsR1oYFPbbc0BBLnHTkvxjcud+L9QAwMh5h5215pZ7I+XU5ScTu55Yt/jwav+
nHAhoNy6M/ymw4xdWgzllS0x8rmyv6z8VmdKsnHXitjh1Bpxwdb8Mj9+FscUTnx7
M0lk88pc6MMh6Wc2d6dqwn0QIRh07bgWt4juuxRHEaevj/ah+xHlEl8JEN/69Cnc
pSh9r3hLt4BZmDolmeeArKdM1MDFX+4k/irdFbVx/7LdXsTpSBcSphMaWk9rgKXz
QfRg4mMveAYOfw1ehHD8GJFYMXQMR0u6hHpbbaJPF/sJaymT1lpDyYhF1q0sZMax
7EvqS53sJo6RcYJcjzX8YYnHBGQ8LWyaoFkCr1NC+GZD5Vq3h2oR74+j2BqUyuHx
ycDpcC5dBRhEST9wvqfeX1uOMs0gcSA9UQrTcMr5r7ddPl+S082KbgRKaXWd8lSg
xzhcN7sE7RbTNPkwHSl2SgsXRRLtEzI2QW0vORj9q6ehb1NX1Z2fz7UllSGr05Or
JNgURHy28Nwg6WflfAxk/hXMg3RlrtN42RAsaUJrqiKf5bhFUqXHZkWKZnL4NV70
dy68gnFJ2tkAAaXs072Um0rADJFI0HJPzeqW4Lgj8QF0/fbhjcVWMBd4wU4PQE7d
JRHqxYeGlK7Nscj6TvosTa5b4M1AtcfwD3H6VLi9yYoU2XImmiTB7x9o/j2HpPDi
T8/eTm2ugXjIbwmPsaPprxzHUw7/+vlNIl0kMv111/Wh/G95f9cwisOvVq8fHv+m
g0BQi1YuTzyxCrDx6VMJ+BrXKdHkupOTKrH7AYzftCgot4LE90YN9ZqL+q69gILl
JS6IaHJPA4W7ymQot6GFjGorHi5BjrY2b0lOKtQpHy0nEoRrI5t8LT8VJyn0UQP6
AYr2Lo20n+NJu6nGU09dChhi7MjT7IWoszAgUHY1R/MILyjJiwjDktTvcrmyA2iy
kg92FXIGtZOKB9SgaOGChN4+1vAWJsCPCGcmIVNdoXx889yxpg/t9QpeaVfPJQGT
I2BHbrtr0J/EeMTNnXcfga8k3yEeE2QgJRgU+1xTwxj5B5m6zm6r0wojOabuWMKc
A1+zFN6m8LRutMRM+mQitNt2YYPKmRd6BUe7JKhpm9leErAXXa6Ob8UIOZk7BxCn
mq0HxNkuzf2ijerHOBeoCFB8NRI9KVLXIdRyWA4C/KZYTHzqsMsrTkDp+Rc9NFo0
tow6RUEPfXGm+FPxODhLPDkmzlOsVPTZm5GOhKb13m44GgSP7H9/iXF0k5anqnk+
h7tImAzrXB8dT9ULhw8HiS1MPaHuLhA8OyMGscZAhxVh3hqqPBxOuVnoxC5rMUaU
JAZzIAYKg6/HG849LLS2hqTHCOdjzWeaOeCtxT7qRHH8ebYlTj0JD/smVJxPdaAB
TWTqVQRheB3oGlQq2aAoCN4CgEamTen/Ow23lMb9I/ac+3smqTyeeJ8JEwqxtIGZ
MMXgAm2QfPulByD38vf06u8vIMDPXaNHcfRELXsT2yOUGr5NXH8aOqNc8K+jarkS
wKsykfhh90BdTOzAbv8sG8YBFYsNKo7r4wgt/9v5QP58Mii5ChfJbXQ/BylxaA3h
mFkpFL3j0Fe9XsM3Yze9zRKlu5JJitctcXxOvtIsSrffzl9xIX5NpUwYPAJzw3dx
TF1LY+oDipRjEkM28S4mpBXK87bbc7ieMSdRenuR64jN7Epr/+ddal4zsudmnOM4
fzHHcsTF/Ra/MtSeFkI8idZis2o0jAupbLyYynzgz1Frrff1xpQnqOwBwC3V4KYB
jmG8jWoa+5qB+BmAlL98nnw1PD4sYg1EBGO4PrOaGRHTRe0AW9MpjSnYsshHJoxy
MFVlIhSzhj+e8mivs/0E4JveHRR8caSM2fBqfN7uhvoLeRxDq5x3QDM2tB3u8otG
+rG1SS48hkIYFUggJ/FQeHe0f2Yudkh6omfMgyl+dpcIyAOHSClpIz7zGrF01VJv
tX5tx0DeGi2RGemUg7QM02YB3H2DyQR/RpgkEmEKIuatzyjfFAa2nIh/Aaj7lnzT
4ZwPTWK5bYAOYT0TBjLKqecyCjYy7qGbe7SgG7fn1Iyyr6JczmPdycq+O50aUJf2
7JRHt/mUfVHA3Sw2+WM+L+Oy/dsZK+XgyC/uMfFyXtR29ZhKyNgFozrAygkZEn4W
0eaUh9EZxtEcbF1fCib3GzqCG5GGqc0MtYEPsNXv7Cx7o2KOEaImayFccb63N1rq
4KjRz5MTOGfCMKSnBI7SJjv9/pqy1VuWkbA2KEfOjv7QvSXkNHZCgfYcMsN4M/Xu
pywbn2QW/VFiHaE7Q7H66jApK6wJ2Ox5PSFhyr+ri4f3m+bN+mEPU6lclPiavVBL
dx/VlxM08xO+CETzYY9KjyyDn4ZqejQhW/wwL18rHwU2bg+NtOiw0qVVsmZPcNfV
vbxs6Z8x6rmvk2KPd3vcDD1sGU3CL063ElOTuUPcq3xKiqpOOHUx0lemyzFnMKX/
oNZ7CLWo8+nKzqg0HBp/QansKBDUyCpiyzAvWU2cfwe3z9RqdAsxQ06aQSWB8ffd
w3fhOEMuBfvXKmU4JfDZJfmyc6foGldtPC674YZuRoUg81q+rTf++vRl08Pw1jsH
u0tg4rVn2nISMoeDka7xweIJbpAuE5NX91bkbdRwwkZIl0iVa4v3KR9pr1fJUpfL
PFZUTnCH8PdR0zo5xPrPpVAAwsLJDRrSlnaFmrE6SOoYWgZmZc5C/eySOnAPHO3g
RlR3r8snHdKUh2pK+WpnEjUFbBZpu/OXWv3QTJGrBMYroyGOGBgJLLX186GiMTSA
7W6uleS9F/mvbmvgD3PIeUYcT31Mm5g1GPJdzjbLSnSiKyUZXyiD2CXk99w1bCAm
Co4xstSp9aNnB9nx7u63ppBpUdyAaZpD5jEwHlq/3YvR3ffvlhT0q8AkC4GWGL9G
B9ZuShW0FVZwIbHh0lnUM3IPG+r22X/n/QaZFjtXzpeTR/+LHs5DANPBo9xl03Tv
sLwnxIkuMo2Wxr8QPSd7C5m6YdmUMot6nTjeLy8027UuBAGX/JSn0A5uFUXGMzQx
2o6diupOuXmJd7rXnuLC67Kq8MT63ALOO9ilqn6VlmDcblq0tir7GAayC1keoSfZ
cb+altySkJugrw4VlSSXpf7bcB8ZwXGs4744Ag/ok6ZNO+vzLH5gNFaFQY0CLVEB
+8nG53UAqUu2/aSHkyQ4JBrMSFi67+oo15AzDQz5Gr9xW6mUwFyUFsPqugeVKXE4
3LMokrHcJ1OYc/THxjwZRSw6wQlw1igzkpW8egCT1lEV0wy/gHyvAntyMEqSTfrj
QABX6E01zXd2xNRVgQC4+PjFX8Jr/15RBJbC2b+M9FWIvwL9g2PpcE+VmksRjbD9
Sd4T49q0zuYfdMyxS8j/G39wCMbtDsq8kwZgHThOVF4hYk4rZmcBCQzVVuF1Pmol
+jln13WU+u7zJHuk/MmbjH5PbeynP1Z3gA2T2H7ys9joTrO8q9GszbEiveCDu1g0
Ro9g7N4wQK2NasZ0lRmNyLr1G8RKHG+ujTMNVP+D+pVeu4vZzz77kxy7MwWfzY3I
pGH8BrE2rZWlU2rr7th06uA/ZVcl87kdo7nqxCp0vhbnk95bMCnHiw5CgvvHH+ei
yYsqX6v6aasz6TD2f3+dyB6V5gqblIyUFUViOP+yqjLH9YRe0+FueivgxkmKwZT9
Bbe1rFs1QomccHWvB0CXKtL5iYXmrv2/kX7mGc3AeFFm2k2qW7YhxJzs7OHGjVoM
z2mmTk0QM8zbsL/mbdX+oItSlyznRDDVomR/pBjTrF3ErCtUwjj5YvoZQLZa8NBh
nDeZF0f15EBF7m3FSKYL+MoBHboj7HGfWFwCkWbbCsFw5/MCvdHlezCs0OpjD4ur
MmST2iKGSpl085BQNnLIZfjKKHD/VhvNpEBp2ms4r6o/oeejvic1bscwuf4t46H0
59uhYpUbwrrMr4gX2+pYoo+xalFZaOqFHw5s3fZGU5jO/4oR54Q1unQ8qNkgG9JO
t7A8Ijv+jr+BTYNL1Q6ncAatZi7MDu2tmPnXpcvAUAE39WSFkg2kQKvCQ9JQh66U
vn4+c8IoMI44HzKkk24S6cbasC5eKQmDGUNuqdn1UBZ4Agg123L04g/nqRXZgMmW
RA+us54PwcwLeauy2YmizrsLfG+7tRzo/7trm72gkX5TvKnmDGImPOGJOaemm+0h
93delk4pUShvT62KYmTgUdA6Nu7s1BlBIG/kGIc5V+OphMiTecYDszkrVPVmI6AB
Fvqrlj7FivUD2NDDlD9uWSrLEd1TJ+3sYzzUV/IyBJSrFT8jU4KeYm7yT3FuY6Ur
1vqxgGklwYcQjIFJ56HRccgycvhDjLvszYSDd+I28EkKDt397aF97QEnVZ8o2WVt
cQy7ja182OUmCm+ZUU3k2sSWzWo79PmsX63qGOyQVwYUL+lPgrWzW6Pg4FEMlX1M
eGMZs3YzQb1hMhCx5Nwp7fHzrz75Trz/KXiYD/8w+ewrpB2fElQbgNY+knVLnEzk
nEdCdF7UvSgOJ3s+VKuWdEeOXXYU5s09ASyb8RfLdfBpNFydyBFAVcv5LX/hWcu9
zE6YwRtQADAP7OMcS+DdUl/0dhTXn1rmWBCOKRbcR9FKZCDfj8vu8Fqu9mDZcYNM
tEGeOyJu/CTJSTAVktE8bwnMKdCVxCurKVAWJ9Z4p5DK8o5MqL2JQiDXqbhHS6Ym
8Iihadnh5OJwAEbsPROfANbrcHi7AA0wslxDs0/Z1JoyL9Qw6c8tnt1UVGjUFj8U
+w5Jv2to6yJwP/QEtOnZjo/vDi6CVJXKh3hndrIuk89EnCyWUQX4HF5CnHNrX0J5
R0uZ4Hx8g+a2dQ2EilxHPPrPZvh5l6aeHunBxcn+aAs7C4tlzyfSUVq7UmsiCCjF
9mHqa9PnVpam7KMzEIYq5V+qK26hMGoIEDnmtk4azpZ8quVl45NFqmMIthWTEiry
/fnpDt4f+ne+LOBE4Df4W44fzxfPO16hK+LLxDKDdTzVVQEsgF+SxFHtOMTBnVFj
iwdOi0TuDBw7jIXzgvzR2SPu9BIvOpTyUDCcrxoGu04d0HhT9AkEJErs3oBR7Gi7
cDHyaqWKQbtkIIsF/84LHLfJoDWVq3LPo/XG22iQQ3cKTmnuu7zXdGbqOp/q2pUD
mvQ57EB7MyTT42XaLXw5Ayq7VkbFe08fT9c9d4TrgjvNQ5lYwrEADg/rYsOiItGu
q8rK8LeHUyT573og0TdWOAo209tFAreVZdpfMaCVZnyUTwaMEp3Q3V9kXWmSXn0C
lfIIQUev8FmSK0+IDJ+WWzLEnY6Q3wI4buwFAgG3xb5PdyfA/4oUFUpEE7t4gl/B
QRhTnHdIII7qdeiR5QxApTEJ0n8EnK8UN/5XQgockGv/LGXzYWBvNtmkRKPaTnxH
SsDoQ3bDRMdDqomvw4xO2jWwdcARhZqrB7nIk+0lbiftj408R0u4VBdL+P5bBiT6
QLgpiG+rwUo4pWejBFG0yktjatgD61/tO/VeO45oT6V2F/gD3t+k6KcVZRcH3uWz
OwWCkEmGJ9ByvVddQjdvASKSbfmvoQ4mS9WsAgxNzldh3qTaXOgjCKa93IjzSCuf
S/n7ICg5mXPESjpSZw6ylK/4XrfKR+mvZfn1GyOnAYTosjk60G/2HAAlAsi8cKw7
7zbuIuZY+a+LuN9CURYlTChHMXh39kQQYhePAvd97QvP9ZOSjv4fc3qtb1TMeZRu
seq7jC1+L3av3fJ4PX420eyuFl4HqXohLDXEFgulxo57Ta0XSIT7wXZ7DBXcB+Qj
NS1wnlsvEBaev0U+gMRlI+Tbjj1uZVV7oTgmOg7Opn6VxYptqtpadddZd/I/9Aog
qrVCykaIrzSRo2x5lZU5eqg8136jSpIbU6Q60vV6MVZMmCUuXV9TCFgu7CyDz7im
X60po0UPqNhTQqzhf+ueS+4XAw5iK/Z8z/DOZM4tBG9Fr02ZiTLPpDyQIFcPqDaF
4U7liCHyf2ptTm+F+t1WQjyfiWLrdooA/F1D4CxhZjq4M/fUEVbK5RcJpxTXFqvB
9hKwWEv4zivYpUe+A+SPsq9KUN2isDgYqm42mobgaIqEY5x+wo9diR71EmOrFPGa
W6MLwt7M48ySDp6ysPLAEXdeDc5pHr6b8u8QKKFG1kFolVp7EPfKtKF8Vx3FIkrD
6B3yOnQJuhjJMG3KK19S0yk0b2IKwVt/tWVvN4+lq/nY9sh1VbGdib5AeRmIzMX1
BXmwC0j2M7TdsRczb3xBr/yG0+Pv+UhK7sZqY80CqVQbQhWwEwE1UFi/gWenFkUA
OEWixtrXPhjcd1h5RF64ngNvWdQpCfbHXSpCK3oWqDoBuiu39a6y8nY3fNLJ1clB
pLPxyXcXObQc5Y8RcVCldmb1Yk4b/RhNhjeKIkYPWlANVzkPlg6TXSrKPdfj4jNM
gpjq/m3wMzerVi8FMrYz3XTc34iBauAs7DMuEtgMduREleWvsPFtXJvkgfZvzzop
WaNkwm6fnuOdIMNxmzlNo//GLtf9AwPgVhvk+D2R7mHbgeSGL0f+eMd+BcNSrmRu
ctcfRr7PR9MjXC5mZgLX4h7PSb9tZp6uaZ6i/o3KP6lr9O8WYuntbp3P+0n+rWAa
ewNE7vQgf4OIr7SKw5QTPA2MTsku1YbH6NJwOM0nxKl7xwU+6gSweEuLTMd2k/Di
9LGRgo+7Ka4oq83MNTj/L4Zt9AdM1fcMTl/hlPL/nT3S/LnySTA+4kd+NrMV5/gY
g4mZaXNPrLQGI2pjB+M3AVO1nxfr4dJsAQyl6jgBTnVv4lnbSTwIpYhqnf6Ylqj/
S6XM63CgRM+IPZDSQUiLGrK48UYWr6ruDxD9ia7cqsMg1zdVO4mXE757hf9szEjf
EVNUjBPQTy9ONcB0/n1+LJ/CB7Cw8tmSNvHCtjpdM2QcoL8fSJUFQRVe1hX051I+
w+kMJeqvxcJEERos7eHUhwbWUAxs4xlja8QqFMdkKkqL0nO1xok/pIN6Th1MddUc
q7sX/Jt5Zf44Rt2grucJU+/a4UeYuyKG1OMWdLJmGwYtS7wQA86xgHsh8+YWaIMr
ji/WjgOthpZl8xb5TJJhCzg9sJuy8YtyxGyDx+vXDZZL/7zf2i8WtR87m0+QZPa8
mStWIRSfI9p1uLSML7TlhRfnKlvuodE29M2pRebv7/iZ43pkfNO5HJTy5GNvxVqj
HIJxqiwquRflKSGGO3ZuG2pHMenWpNR3USbdkJmpjAWfOfjGFz31N8psBsxrUcMb
CzTLZhImyH65abuK0HRlyzf3S2BLMoDVkydX6E7eZ5zC2Q5l8lbUIlVWTrBV/hZS
udtWViyfR6zEOM5GEUcpwvgquF5HMWkPGYhGMQQLVoIufIYTP2vUwutW9PxgF8H4
HUykymIaEU8SyKXh9ZW7QiCdihz7RadhIEXexrfr/kGY0Bt0IKCbc4ox2KiCkT3a
DVv0b+1FaYFPWwGe8eCvspUb2ZNRHVvUSLqE7zC9PGIkUZ+SEnaowEfCgmTcGEFG
k0uUsKHfriKwVdJvJrRmQqCvtW/MgHGQR7tLzNnFcmMq6yiJ2vXioIA7Dw9n33qF
Ui7oUks2jTxa8R4l4n9fsJXu+NngnHRBC+JfM1lj/M9uBR/hmD1vqspE+HYQKUZO
7pDF6cEUwyTvq1kpkEAtw9W26tsYFk8vLn/nlArCQZ4N7S64QF4Z+kr3Zh3YhmRz
Ktg9N3WllawijQlq/m35gL4Uts9Dyyz8OLBkgW5579/BFBrY4R1cJlNQ8yaRD5QW
sk6XWUqOBw0hgIsa6Vcjgi7X0LR8ag/Jds66kI5QTVh9ATWE1eScPpI/CVOMkVnm
FEcAFkOvthbXQ5hgQUIyAfguBNOC4AgleTyItRvFCVVvsyfRRGCOiCt2jIjAYtqT
nwRqdQE+77XZwzRNvP0GgUNcOrSLBNqqrL5R3wl4Nwd1vyeIMd3uyuloLumkEN+i
c6BqCqWdSruEpNw6h7odJ9LQppDHh+t3qSFHbt/C84hI8cFWEq3vvup5mIASKry8
emsy0GSndp8dyetIKM6q91CgPcw/3nsSXFbC5gdrGhYJDiQAraVRyl41drY5bho1
ot6WttVNqzP326gMBwrzxflMsuWZdCQI8uFy7/DqPgmVX8dispgHjltH3ySbjlGf
4SYpKk+BIHBMSBtMatkTqv7nQOlZVTBY9rB1OZMaSo5J5pcZXlpv+COYrPVHQB0A
I4otEwAyVnjjjoi4R7SNfGyOxVMqMgt4mq2ipeVeobcjJbho2RbKGeijLWZNk8ev
8+upOtd31MoIpcTfo0HVOGUpX556wiztgpb+wx7S0MLS5gWfYoIRlC4n3k59QQ5T
AMcRuHNkFP/D3Mw5euuy5PdSwYunmVCUKaFQ6P5xjqvEkpIX3HfcuUjvtWL+lxXy
5+nf0ks9QhpWLwa9rm+46YHWJkzsUu75F3qHtT+mu5vB+LNS3N5ruN4awa78uWNn
WroEnW8GwyKhsfcxUmyPgKMzGOJxawWbEVdnTrK2cgvCrg1rCRiXf/54CN7lgpc/
8Oowg1nqxboRRRaHszGBvgWk9spFdsQJ2TrH7A1gIW1vTpsJJxpuSlIoWNPuaDU9
Mr+9E6Ep7fWgHxaPO3kLJH2cxOhZWpHPjbhf7p9ZahswTBofS3Vn+jkJZMw4ffAS
9NLSshgRtkpXDXP0X122TygPF+VLvCGV0pvm0wgSIQL/D7no26tEOBc6GwR/m97v
rP86PUkNBO+MYUWNaEb8oGPB/b784bvZWTwGs2x5EF5mzb5R5nQbi+ss8B2U0zLG
unWxbLk03o/jqUVaixtlZzto0wvKsTKXzop+dMTNvuyTNGsLbhxskQRhioxGxoC1
Af6MEmOEe/fDard6AVAf7WNn5lTa3TA98lOYlhtGP8o9CIFd7IteRhRUW4yD1GVF
Vh0a2kYms/LTDgBl7zA61Vw8CcjfJA4va7Uzvqi7KZO06LidEQSqHqtAO91Wg3U4
EBl3V2muCduRr4d4Gdrx3pfQZgN7TJ02Be9Aurs+Rv4Dn46G+ufNza2NnQvco7bW
wBmYyhg2pT3qhLpKbrJ9bn06g/1RWDTS/3nT/rouiEGODiU5INKbjbxmYLky+347
9qIpAF07K1MT4Ur/AxQMBWmUgygUh4fR7Q+pSa06rNh7SERwsGo7DXmFiyxT+xtf
N7QON/e3wBR6anFbv2HS0OyccOVc+KNGYq4oALyQAuq8/PHYyC8zHtg6SlmqqEFt
OiC0n/svVRvBIlNmpL8Mu6VgHjE/NhIat5EPyr6Hk4AgodWNRA84EyZxOl5/hScN
wAH7u7wlzy47aEv3xjZ9Sw3a9i/2jo6T5kF5Dwi0szg/xcwmzsiKMg5mHoBQFmdx
3C2SnR0j26ZGz1ZWgZqF0MKSN1WXAauLlZP2N8KetcOiO4liQyzuWcr6UEWPnRUq
TrtZa67UWQf01dk6/0aLpT1bDq1f6ek9Nx54vbpuviEDA2SWAUAkCbvYOsJqXJ/S
p4xq5UKNnLpfzoYAYmrpcUMmANrfeSOphd9cHGCSV+OCMdHfI9nvB+jHD3sFFFY/
GmntTLdC6f8bikn3pAIWcmhTIOtrh3IUgyX6hK/XAYf+ZGAHrifVm8uV96+pV47Z
WmPjwaHPP6pSZFA12cHjsSEyH+Sgafh4oShuvrNTayuhMP9QPyA0gd449whrQKoP
7TfWn/9tkYbpVTLihjomaz9dYnUBWRG/edgURG3MDm/3A9WGd/Exx6G4ICQ5LsFT
pZ//hsZyk5qoZsjaMN2NH0MzOsBGWTwF7jVXO+rg8lVb59am1iecZT2W3b0IlHpD
+moBGf314pKl2kGjvdQT1nP0+TCmSCYsByqX4crj+rge4nHTh/kQWzwqGX26GtwC
hKiH9ptc85L1/QjfjCgI3GHzruixJHKgtT7+T58iiNeKKH7Fj9EFoQgWr3l3yqfg
BfpaWZW2WejlmJCGB89VBAL6Hge6qAFwn8JODybdrjayFmSVDiiBQ6+NzmYYSsFO
RMIHx8dJxH2eozbTcJaKvm7OQwYrzcekGr4GfSxttK/GfEkFyq4f9fb6wAsUJ5Nk
3kcdIZCPZGVHZbo1SWPMVQ/JhmlApfyZBIRLqWRSHHDr4qh+xFbf35fRXYXwOppj
JFyBatZMHgRgAFc9JIBTudRT6x9ukF3p6WXf4CzfpA+juA9/l+WDipKFUTMeC29e
ojvIWPg8GSAYg8PDAugNFDQ11L/1OBXi3dCFre8hesjGxir4zv11OU1Hulbs9ZkM
5H3nkcmaxuW7COQngMFhOpdMuNuY99tWwnkzuSfLYRFJZkjeFmOwe0yS1yRqsXj+
bWrl/jT6sLvDOdbC/Clx2d1ffqAT7S/K894/3PxcbEvBUEDkSlSy5TpFj9Y2AzLr
PSGUahWevN6uj321mjeVMUNgZ+5JulVLp+5kmMP5Kw1UOvx54/YUX8jjqR2hXwN2
8hSKpF7GO33n+TTRZ2q+5crnM2uPCviWWBLhIMtaW+xcxtv8dIAbnSbIuSJUDVr3
wRfGaIl7zi/gsatGc0LXJ4JJahkU/6AYpVhTHdK6lsebrles02+NBlhFPwWnMb7T
0jvqHPdQrYIzwws2vRCdVK7EBaJ7WsfeZxR2FN9VafDCchrROxGZWHBexXInoibB
LLgsz4zIO4bYuQrlphQhAevE+re+zG9uD+0wYSobZSE1f3oWypA7SvG5woQzcZ5y
lRA9EHxelAo/rD89asYqtNibllIiorYgrRlXFu6WpP4fDFJNCzLnR1hM/vAsyWXZ
7HmsagHBJjBSWVk4dDSzeTCdufvjFEhIHecH+iDxctDB/XJxWYpniMfNWqecGtNi
N3A5rhgMff6GJsCCIiErslxZz3QB0oGM9w/Wl716lYt1YMzTo+LRV5+xCUAyzbeN
t0wPjJ+Qs7a1kpy6k68KDXw8hW815PVNCJy61QMDQYWl20NLrc16BR09Eg2zWBi8
YqglxzaDAVtUw6YF2vrd/EYjSSY+O/z0UMMkq8Kzyz6RgsBRaIIdPusiH9VLj5oY
IlyOJr2MiTfGDb29PlDoqzoo7niKoNnjyDxu0U7PTIB34zqzWlXEssMizlyGSqf1
tQmPauK3yk/fiy9O9PBUgVWzTTGUtjQ7TOHg/F7byWsgf4i54mkc76EZIroegHTG
kkLMPpvkUFgnu26mQJzvF8rFgQjq2QJV4PYVyEsLnrx3kuZmWwAhhyDBev5zpUbw
5pYzRU7oEZK3mP9r+cHPJUEAzZOOgvBcpFFFWxG2miyM/zsc4SVJZjYUy3P38r1H
4+JbFau9cwrscFtpFxnkUzG4lgFlOT05kEfcZjM8QE27szrTfGBJy7kMT4C5cGES
AZzOvYF5ePfvrjnPnN+iF63vASPhXpT0/6CTa2BPKXP6n3L27+gItCMufhKLK3rx
29/yV76FGgjs6S67AMKoRR7TtNCLTrjIy4YMVePb17ds1E+tpy4pyHSUdoGnL5Km
y52arWARJvroGd/3ogEc3mYQvjiYiV87+cIO32CzT2wJOWh2YnbZbL7PLuIZGJBi
2sxRx9CeP3qo+bYOXr+1oIJ6I1wD/C5bnvhvZNRQJM0Um5ubwFAWAzWBrLOqALa0
5hWtFUNxBWREIUCJiP8lr+yic9XE++l5FEmGbByTBQK2AtVtGltE6FgadKqQj4jr
n/+LXG3YS3snqOtFwIXr0msiVuGpY4wuZY1SEnwmk47RtVqP8SswAV4ZRDnrzKcm
cg1OempmuUWAbKNKY8ihuxvA9p2jxL1DSga14ij6bWoR2yblqJvHtoWThIxw1mYg
QqPDhlT2zUlmBw2C2Nu3TAKYjqILrbRNyk122r+s+OOSomydNAY5tMwmEy3iFa9E
8zHa0fT+TfJPq+fXKIw2hYBLw45Y47x69VNdtQwSY/iIDGIRizWGJbSlXDEBT3yz
wizUzjvquX0AGBo26/Il1Dlmoq4n6ZnGcenlWSwIKwfEEsXB+FN91LKtxbgaUgOm
hT/3Z6svBlVUPHf4J5h+gC+z4+DTYiofMXQ3nETAkQfuci6h7Yc243tFVSMOm1Ah
wDtCqYY8pm1r9xLhH5fcia5ICW/gFlplTNbqmBVaBghz3t6C5wPH4izbvpUOml+y
m6ukMMH76jIQ4Ebq0XsoveK4Tt651pxW0KieQRxEfBoj56mqp/qnXqGheGKhiLMo
J/LqyL5Ma5nIL0Q2WkF8z093e5q/NnNGlSChnqrLqMmyePFmcROyW0accVqU+TMo
167FnYkEkcd5kFWJ86Z0ixIjKqlbuG3x8Vg88Q33xMpxOFPmwefBxFvpnhctH0EA
XAIEIOjdbm2/ZuECaLMumRNngXsLO9GjdfBxJhfoWGnx+w5ykgQv1n/16r5PM78d
sHUfe4XdFI0tQhTDgA2argqzteZkMbR/INB4GDAEvdXWX6HVXo0NciwDZWk0Ferq
QvWEVcU1lPj+9jGx+uPVx2KJYGEYjdpyOqa/Grzu7FyFMSawnM8Sx4UIcTW3BCzR
nwEbXUSI1mMf95y14GP3ChGI9sKwKfuO4bIJ1DWVwDbmZzjjEnqlBxxpcHYrJKXy
8XHXLDsHcnCUjNCZJ8dsn+x6KBTF3Fa/7g8QlfWgRVvBddEui+Dyok4YFBF468wQ
rBr752avrIL4qw4hHyXm4BKhcEuNapkN6UZ+FjzR8BZ38qIxpW+TcxZ7tySbzG6P
Vp/uyFB5Sr3QpbMZS02x5FhtjUVnKecb6c+C3+0g82PmMyIt1WxipErdOk/KJy55
KhVhfhzSEFP8lx248S91tY1L5qKIeDdl0Uyy0kqdmZWD5uaSNMeMusEZIQ839IU4
SbWOyQFYKnAIZl2pWJSo+blmfGxyYnFYcWEx1w9UpG2ebrILuEawet7iAFzVdfbS
E6IwkyGd5NpfIcQFvrwIPJ0vp70VvbaqTjxk0A+Q9wWxODarg/y8InprTsUMmycM
yt6Sjj2FtTjnEYltP12PP9cnTxl0VH0Yd4/0pxLtklshKeX85OcGgQf94VMCL8Hg
Us0lbmOkfKBUldmJ9VLw9XHBj9jBiCQm5acKCuMuLJqknh5iBM5TIQ2nMmqWX59p
wWfnfVeHdxwz1tEq5yZC++qJKEtrkmOt7ECARw5TAjgeui/9fHl03DU3Ozec60nh
Uu5e5YzrM1nQCnrnvIUqi0YqJDP+FHoMPRrXeSn8S4bqRsAew9BsOIhxTz2fOmv7
lcOFF8mHd2vpepMq/WjdJ3dnYUa6oWTYRe3WeIYlRvXpEkxsuTXKNJvEq7OK2V37
4x1d6G5QqqH1cIS+0bXIWJHaaqBZhHFh25CPWX8vMh12WAhvzgP8vHVdsBnpaD9m
BwMPugMlaO+L3bzPGvXDdUuNEpwHZpTP8rYDFwoWzKRsSFjzzaQlr+9cR8BtO8cw
vk1f5aRDp2QEqBnQOn8Rj8IL6mm9WeKX7NtHX+SmkFYPIavFc21U958oIqCOnPiz
wzqt2iESEHEay5kejSeZmNO3drvTrwr68OwU08VpdV9mTMAertuX8BtiueDEVFyM
vzpssajVpU/ehPveCEHFi7L6HeNNAZ6EkJimfcq+NT4q189CZjRDPQD40ODZ4kp/
4xifl7nvHP6iPfJuFLPyIto+sqJRf/Olkj5OkmZCJ5rjlMcVDR8cQy7pvY8lIYig
XHMrb8gUnf3LZhY89ChfNqJjs72VG2WN5PV3lI2Lkf2t2D2w9m7lnvgUf8C/qJux
VYNyY4G7qguFNXsmpNGdy+XXJs0NS9UyaSFCaeGCDEuwcw1a+MEVPi7PNTcX3ovm
5cFlQxxbPO9jdFflh6C9iRTMFcvCNWRUfSpXJRpjAKyKBJFBD58UCAnqNil9nvkp
V6hnm1Kk207AsNMNMBtThq8L3DaIFN5iijac7+AShDWqAt+2HfXtRjJ4WH2jBgTc
KyxfgG7NvHCIks7SmudHGqHcc20D53m7/9uXFQJDcyHOni9Z9MzPufj/IwTBDeGM
JbFaApq9RBeerVDmWZqUdaOnSIJonotTx4t5GUMW8TMj8ReQ9zRtvNRuTl4Wte9f
6NXARpNja6wcR8sFqrDLMZZAoo4V2gu25Pb+anWojZDZZyfsIs24TRJZc3k2glnN
vw/wI9KfWYKLCwdZV6bZzmVoOy/qMoWThwXOpOYOnRRnAnKcjsSTbBi/EjZhMNmT
qbo4VqHOAF5PD5CrZFJZ2dRUO2iapjFeAosr6YsWC5Q33Xf7XbQERF0s83ZCgSIb
CzbN/YtnhYWGPTBFiAUr8NdRrqXlZDkphfaFlEwWyweRKtPbzHSRn03kxSkA63Cp
G29YqC7pT2xdHIVy6hxrFA6mPXjYBr80AE94w9/o798PSs+AfBtlhZGbMhh8KzCQ
qGmF+bssiBtIUx69TvduF1ssXLbkpmvmxUHPxQGWfqCAuNaegMkvi8H4Dop5emmD
RyvTWiuUMSxQ+oIamTGAoH5LebVc0UFSUONeROQMd6Wl1xbQW9x5ktcPWKGlet6S
KBIJQJ1bpKxpA/bAf6cMiRUVS9iL78w+jip8bPhbaY+9xkAJsR64oK9NsSuQhwqL
gm32Ia0zQx6MVQMGNxqRKyaDMB2O37z7xEw5TJueaoXJ+3KqPfb8Pfk9QEsXkFle
wqph8ICUl6iMTDPit8BtNPqNW5Xqf4bbqpS6Ce4wSlCUmtELfDjLvo6+OkcRDtpx
78cfgsusrn3MFaEo1woakVjk/6M3xCAhRk+4JsR3YHAdLtR4hJmjamUaA7VaATzk
Lxq1y3DvrGiTNVOO7kWef8gRC/qdqsxFq1nqhunA7KtTuEsztAEEhiOnEAxR93m7
U8tneBeqPu7uJRBHlkJVfXH7AOqXqY7oD7W5aXiHqsVhQQdb+h2mzFUf8StrJgNL
a8l3JEsNNcJLMzDGZ1TgIYQoucNadqYo4zt6VgMGhbat85W1Sq2vpFcFBw1R+iq0
XJNFqoNDbw2Xl2kcVzl8HD1LMsEVK1g/fExafcsIrhKSH6W04HQp68Rn+PwIrvXx
CCgjVX8pLiiFgbwsvM8CzKUL5Ufaa+8jr3OnIJk0q5NvKf42uvYWq2gMF8miNNig
B/ZxVcGETd0kX3/PvNHKCyazTsiAfL/oI4MSPZMxMYprTnAxjURCo7Oxmjp3v44F
YDIk/JdVswxnfkppodHJRAkDUQVYKHQdu2/2uA7i4qMUq84xRdltfY94E1cMZFM1
ZYGMaQB3nt1m2wWoR9d4ZSd7Y+PWTz0rSy/AeYNN+9eHAdauxjNSMDUqcPwTywwV
XSFLcTUDwWUd+4T8iey4cVq42Ic865YGgX7dWWz6iCd4MzjY4z9aaOxvuJRZXs+6
EXSYFaiLyEndxmEaLbAZJuAGyhcgXUG7jUyjW/lBYR1shyIZioYqUm2tQLkKcW4g
iDILfv1Q3dYNc7WZTmTLso/XUOQiLbL+3AJDty65hHYukgQB38L8TkYedu0aigze
Qg5FD3qHg+n/L0UI774oD1vtiquofEIfH69gt+xa7U6qIo5F9t6sVyqJ7emi38Zh
FfHwDOt/w0RfF1fNFwNsRcBmG0Wm/mroYMbjv2QjPXMPeAdrhhC2CanoLBjBOLc7
nYQb/fO3JkM3C8qzpEJ/D3D9K/BOZxe5koSiSsWlz9O9PUOAnZ5mBvSP0j9oHv5O
X8dHsH/uK2V30Q8F9Lf+BPEctVCNIs3r89ryJcydzsFQkyBEToLheZ6YbmN8Iw6y
jtG8W0+Aybjfxs5yAMKSDgsxc/QExzaiYo4HSykcyijxEWhEPLBcmzAxxUiaqyVA
oMm7XlaYezGgSvXtFGrZMIe3fE1XuEFjhE0MD4XgbzkGMtrenOIiMRHPQ8vAbX6T
PXhFBY8RP0FaPSwb44u5u0ZVM8eTF7sC6zkPz+jbN6ezxpxXS4Z6ehbLpR0Lo6DU
loKiIOyundPoXbydo0GnA9eoj73w3sd99KC5GXkxqq/VDhehqhjADM7njPET5K9B
i/ptNKrL6lBBXsdfnVhcI9CKBjn4iYMIg9s8BK6RCUVi6s/GOVYeS7PmNKWC0y0k
wuGNFehVx302C5AwYgqm1qCBDcXq4fKPwpqPwmC4iLIXNNje36ePqaWiizsY2GxG
6vaddu9Z/rGKkH6dAXWuly2HMl3o39ov1NHfonq7iqzIAfxEijOP1uS6zKzqf3bp
NU6u74WJeCBGkUr82xgJ4PHr6hdGJSFg/a6+JtojW97Xhb3yzVRdodV4fq3GYVdd
6OqEEhw4QtxGJVJpyj9QWdloLLYYKsrJWcYD9v1j0ua5Exkai74myccYkXJ2CdAJ
W/8j7vhxYGCgi0aqNyr8BNifANUjkF7E/2R4C/3NzSxn72PXlXc89/3Fe/5tZhn7
dzLrNpOPCBO6l7uuBPvuVjrcrJyAIbt5rsRarrfPHWvmpIPvEYMl1owgdvOmkflp
PrYeaMr+M/rtHnY81liFcVDbiw18SP5QIkw88OB4nH5tTyM47DvCNVuyXO2Um9vA
EGzSRwijrvcChpsNq7rvgzgx62eHZxmZMYe4VXubd06FZeZgO29kwoVw6IHl9hD3
Pvqjuz7t+Gsn/GfW6G3azw4lpplMorOojvJHf6ev5sBH6QCJC9Xe4q9N578M8V+d
0gM62ROmJEEA2ySibDSi928OF1UJFt7Vj2JbyRrKBLk5iuxQg8COiuFb/ecEOTi1
b4ae9tCdie3KsUm96d0lOq7ufTfjTN/0mISqyEivpev1kF21+bGfzeUffqph2vGa
vb8ugU33GmgMFZm3DyEgT9MAZ00sOFWoe+w/rqRCz12jVrtXkLFfwdF2FzfgW5RW
t50Sr0eAvpMBrpJlZp4xdIe4hSPEhIPKlE+AgtLvFiWnTr2UrRHpIGaA3BZtrJbQ
VeD2+J3qtgDg5eJLqDKpt1JDHMOtzIPKm5TLbou9k1bRlTXopiO+m37fcITEz8Cs
IzX6SuSfbazpQ/Jm/EhnFqbxo5HE6nmQ3iJXmOM2qTmmyTg+NRJLT2xBLk8rJSPV
RmdS7AzDoI5en1F3xuS/enNvw8h2ELv0r7iRwmf+UzBgN8i6YqrS1cJPZkaHJxxA
1ozxy6ZH9ol24PVSbEsXXeFjjnb4x6hoNNdcus9wCFOm/Ge1UohZ46pojm99W7qs
MXRk3UmR2wDTqj/W+iWB3hEGpS3Rs2vYiKLBIXxEdKO4NRQhN/b288j2bEwgc94X
DbKOZZetOJq2vtgDQD3wMJG6QC9YD54Hh/ev9aet0qMjdJ8X/MpVRQAy8yVUgtkl
0JzCMLiFU59WQLRfD4qmYStbGu3bstS2xU1NfTSNZDasPWYo5CI5z7B2UHtJ8r/F
L4t6BYepvI9EBqE5A4ZKpArpjgVYeAaP1NXWEGoqe98HJ2I9kcn/C8Pn4y+UHTW9
4zO7m+GjG/DwsntK9/Ohk0H1ARol6lrNR6KT3NJ4tgGjAJOFwYRCjPlJYsiUn+XW
G88Ie6urRA0ttEd8kKgk9N1duOJASloxTJM9mQIQ4z41SLU4FpiBpOF2y1w7zol1
q65NARCsi8bHmoAWp2mOnz8HPFEc9XnMcvUvJsy4eudPMFl7ekahyqLrbahp/1Uj
mErSG9FHEYNpZNHH1WoUR9U4zL/w5cKnIUbLR3N0duVv/t81rLvZoDSJEOafqzEQ
lt1R35IHhazGsst4jDJ/01EHoAf6DeeNcjvgT3Rojkdd3b7ymJqoy+0encmV3gln
2KxKU8pRl/FWNUtMldivOzvyysF7qclyGohIqxQh34F7j+mNy+CWklijIUSgFclh
UtjXJsj06n7nNcFI5Wtqng5w8kySf+L3HZLiV9t3TGLgzq8fwK1Dy3c2VU7fgMyA
ahzmQ2TJQZtombQxfQaMjFO58UKoTOfI9HNNRZDvxAalwqYMbcgFHB8eJ1zSO6FA
QgZ/DAnuvDnB9HDaODaRgkuuX/LJK9MOwJ28Q8f/N8v/P+myMfWHIQYao9WNY2zP
MONro6z2fcFE5VM8YQfQhusHEzscBU4CkhJbGtGcqu+yUT5pGilmCZ/J7OjeOV0m
ZzLARxDxTymV3U/bzlytKlGt0wjqWl6DU3vC/wcu3q1wRzmeYwA1JBwIezZyOXea
+WVnmHreCLF6yzZu+hMTZvT2bgnhbph6vLPGjDFLDviwzyDTxALM3LXuRnFp8sX3
4i8xEf5PxD8zO55FVEpfF7vT8QbNMES0AFcQnfkP7E/sJDZumRG0HitZRW/i6rhQ
cvsV+PlkRtOOvvESfDOgLZJ35NYRwdhZXmxh/ZnKDtabWn1kdkk0QHqpg9YHZyO9
iR639p8O6y76gqkF92eZ5kOFSTEzoYbPk07HPjOE3BpPgIY0mv1ZgRkdzDysidCB
bMoHIbym7g8pv12IJ7IB16eMcI+K3R3SYiECemOyZXyRxJVn43jYoh3VumnShE5+
tqXgNS3jAnRk+yO3iQhpTg5R9cvb3IZbrpe2fAdPMRDCoumIhktHHB4L/gUU/QjI
tCcpD7HfTSBr9ULCMZmt214CzB9vMyDFLfc6Dc/mHAC+bpX+1XfY8kWDXhqvFF2B
arpGTnu+tcJ7dyJJTDgb752srP7iOOf/K9NUVB+/cdf+yCWsT//bj1bRgIzyuJIw
80pTZqZ0zF660jBA+jGm96pUeM278ESlEkhdUMnEwlXhMeRszjqfuTOkEALx3FAE
R5dH71s9zlximy7rhtzsGBfjf/bli8bwmqic5/dRUFxg4UqpwcX/wzBEQSQCP92s
BotKjpS5tZyKZStKxPjd26Z4fc45izuTGjNaSDYcVBqiEIyKKqFxP6p0dhAcopWa
GzKiM+fIx67r97GYi+2FXjQ+wa+mW53bypN0RCc6KGtyQafI+b82WgCKrcyeEzYG
Au1pVVe6ux1kGkHu2kLOw03PqjYTy9P7T1YDLfRIo+uUUcmh5tgthzP4ZJpQqvVu
9TFN5ECTzkGSbYORDrTqFTAAp9W0gwJHTKSljZUz6Ox4mnma2BB0kR7UtHZNEBH0
0bBOmWSNRJ64NUBYl0voevbQrgqTeJ+Z35dhUMhCutWfMki56RvEzT65Srxm/GBi
txoofDB8o9uYr6lpNwkFCzaZ/incO7mD1AxDcDMiVqk+NbIFDiTW6MDCnFlc60i0
JeU2g6AfgwvlAVAGrG////YpIiwUMB2QSrb2zHA6zRjOxowQoig0hI9tukSdqlsI
zOfyQ+FZ1ub9pcoaxADJ8fnvVfwXL0wgczJ6MQCnMoIj9SewyL3BQna+cQwzOEX9
oTPxfZvO7vIFWdmH+WrBULwA+XjH0cXEGMSUj+2n91WFtSGsPqOsDVoq58DJo0yy
5Z5y1LI0Kz6S/ckM7UDHcQ6T8wweqvF4C3Rq8qjFHy39az5PsuVZSFNrmiHnLsJF
/eBrkJtkv7oQtJLHzfYBu2HgrmkEarYEDGRrOUEN5DI9NfbQnQvtv+bxABHnQwPF
YTy+cSUY4YvpH6gq2eTisA4hAmEKUx9O94D/s7nuxaitm9GLDGtk8/PiCiKAHknw
jENUTKt1L75kOZ/4SQuUOTgKJ6xQC4Aroancg1t1aq1xgc2F+j5hm6OskgEfDuZ1
W2NqCGwl69MIRCLd7qcrQk1744dPMObLLNqgi4cwD6vI2ftePJFUjQPPRBOFqL2f
SdSGmYFd3YFlTRQKXACU3KLLjWxRiA9D9sqN+yR7PNKfCEDvUOwiBc0sWeeI7GOh
8UYfJH/dvcDYf1yWQTLPpSyPbrJqGcdCrvSLScrWVF00Pj7zdpr6hWenEttMvcG/
BWgjTaKMCZzUrF+BqkaZLUwTf2A/ildmECjKd1bF0f6zKEaMB/xUp/jSE5Pfoijt
4ExAv2ExV/7jCYe2hYqW9rei35atNg6Fv0y3GLqu52hIVLDkj2jf5GWswroCrOCR
3CTYdI7fwIwbHqiqzSMvk6+oFgjz6vkPmt9Z4CAgY80YCSHURdYskS5EofoNibih
o+escjjlHEgAy9mvl2Qn4BJWJI+Dhw3oEoVs8ZJxC1kLKpnBKdlmYcP3HEriWsrd
0O3BbJVvNW6Xz9GZja6XWzBRTpI9wjUDYqJjhMObW0NyUOLlb0B7URSpEM1pObE8
ko6j2M1mUEz/A/QCwu5MECLYKlm/cZdwsrY7wQLmGY1TMMp8sdlazjfOfnikPLeu
2NBRm3lbZayNWiNGQFuwozYLis5me5Dy7+JeKm9m0qM6FItR1d/WpafkqRKdQyi+
LREPwJ43JUKO7T+7NSBKT21DjSO9Hi39PwZHswq/At0nGY5x0go6hOzZ6G76Abap
yw+v2MPL9bJZfrTAF8E2lxn9xjkSyf7ceWEWyLXGjmPBRZBD4Yv3vwRbbNq7q0p5
ilG6NZLRV0T4uQ1c+16Zn7VVRB7w8SJwhLbtPuU0p2dyj/849xicszdW4FVUgAKw
znXuVFy6uFRT85H+NNRaZSfnpigFyjhHKj2+qu2jw+TLEUUyVdvwZQAwatiFhFTS
6xiH6ljuX7SEfg5Vn5k7GbaMe8ru8yN/nS7jOCm+luSwViuEnlcvVL0SHPHp60qU
UsC3+53JQGUlaGAZJrqVaUPJY3tnMWj444XnTudEAs6n1eNAwB6h9MJ5KTnijkso
2nFkrqLXRR1RUGJJkz5La/CvJ9CNHb3D5RAKNn3gkfUVMKFNRlSEuXr5flGfsQ0A
Jy+mJdAj185BwgHGVlD2ms9j9/nkypeGwoNfj/ieakh881jpndz2nBqGCo5S31vV
IEzhr7esrJVIqBKg7ANHvBp5e8agLCHplLjC1fNuxXRgRZQ9C+/G+ikUpRiPxW2s
S/Up+vAK8EhsfbbpdtCi1vEFnyvG6oMowD9gBRPscVPS/xkMItwAdvSYKTR4o6KV
mHymnGOHNIwLLqWEf9DahSzKT/ewT5VTOZ0FydrRy1U3N5i/kEshFArU8vkror0B
gFEMp5z9nFsNgmRxSfBxJYy7w0zaCsDD30eY+PWKIzQOK/zwAR0Rbf6nlZ0t7GUh
2iN6++iUsRS7GK0dpS7T3kxB+o/JXg/uR9rDeKhMF3N/EBTKJSAjMvliBobIO8z/
ZPXxyvnlPi3nDadC4QaC/W6kq9bTbgf3lrD73qvP02N39soVLI7DmzR5C/YNgnwb
Uo3yRj9oODVPrqGBprkLrgIA9O9bjcJE/brYWcBFkN+5nXX6zG3rWsEBWnftzdez
4hk3Wlx4EiIJXfQKEYcRCwhjZHVNWf1E5+vUe+z4kI/STIzPGYfjZXCPH3pqOncL
rcz+nW7a0Sy6JZ7ZSoFqWaukYcMfx8H89DWykir2WrjcKDncRNBSEl+l0UcjkFjL
pI2XciDELhq0F9hxWX8jNaasgOWR4y00m4lXHD5O+K1DpLvUC8wiSrWKIrYECPM7
ZHwsSf+Gm/WQUmjSgQnXIchyFh5CGTLF5Tc9cerZ91LNMT00AaDpQzGbaXQQK4vO
R08N6NzBmnQ07N7Etp/RvdAgeHXELFZ/AG1t0ovos/s6SjjAe+FHlp9QMtx4cNh1
Niniwgh7k/JQexOYsnKxnPINlg+5GBrFn51JhL4br0yqH6VcoJm1bDWqu25dvUY3
sYLxwBoGzqbJAIJ1EDqkV0ewfCBFtWTuQIKsoDogwYWm+Y94Xtfy6Yy9Q06x0TBc
zVIIl27wYGFbJ6fef8xUPTbf8XOApRl7LfXRq8VHZ1X7amPPKy7RFFkyN8KZ8RGz
Sjgx4SXh5r4hGurYvOemMp90DXVvwZZE+KOa3qdnlesAgIbRFhIXUcSnTAqMm2SL
xfLSkKxETEN6GxmPFb2wp1d68ANy2nme7k6vwUvQ+vAcOGW4VKjmsSt0pKn0/XPU
PKFOdpWqaX0wwLe+aOP2IZtmFpEuSB6Lq3AZnlP8XmxojjvnpcNTx8lvWbr3nXA9
ubyncNfvWXcS3hAvPcfgONzHIbbZzLXdapxej82SBNeM7Hfaa2t/VAUwlU1WkuBJ
j6TF2MQAb2tAL83CHmht/VFMfYEhmines7fLRrNX0R4l4gWQenmeV1s7SDonGWjN
uG1dZllvRyM2yCPAaIpzzv0aSuLqP8Czt4tHTL8MTauKLvXS5HG8bEWY8NCnvvE3
o6VdYAfkdxclDp22IEW0oUPOMT0KXb94ie3PwfQyS16KodILdGR0IlnJbQ/muEqR
8dU2fHH1Ws4zwf8FzsXf1YO+OIUB1Irumm50eyr9Z4Q7Zi6uiomH5vyER1uB6PQU
LCsMBaWs/rViz42BCL72t6S3uO9Igu6XwCtPdFVNrwee+xx6xoNPPYQifS/uycPO
34aAg+gL/afWKugDt8zWAchE8Wm1NcxdIhDFiTJ7D35nQZSBhd9T190fx7ap+OvY
RYBa/cOrzfa5q00F51GKYHISqOj0weBL/7cYkyWBbDdmPsS5VV+nGzrdPygsM0Z5
b8BMfmiyVR1BDvv+aD2sVoafCdcUwDYZHIYX6gdbBv6yw0nOlgbXik6M+Q7JslG+
AryOiGTwbAdUElJCr8cg5ZOq3Fhk9+3YL9Ry2H8nhaqKv5Fcw1AOPSlKy93sZJaK
kaGyy0fmJZNhl7TqBBT5zlVQ7CCCNrXXkekGVCx2vTEbZ64iKYEX+/xVCQtWGjty
Xn99uoc40LAEGS57BZHAUf0L5mQFxMuemAijaa6NSekgshLdODVcxiGjfG4n9r7H
LgN1VceEpwm4bmbf/Vsx5gzsvhjxOij/iReVOEuKqBIzvc9YKsv7EcA6mBvQ0Dv/
5fqvwDBRL5LnZry+gElbf2hItGesZVaA4UYtWppkfQ1wJsE6b0BJW6dn5eMChQGY
VpvCYupxgtIP3xD5gL8s/JKvVHMblvuxmEknT98ib1IcMvQNrj07sn7asNegrLdC
JWwPLbirN8BOpyQBfuAeSVZMN/NL7q4HBuJNvv6WI5IjIQGUTkFQsEDw7/zuNLcT
0R+amKdVAllrAJiLTtP1CPvHQvtr642O0VqLop0venpQkHhGxBJVJ2wz0x2fgbYE
eQIYwJaGLqDY2anY96wG98UQhyEifgnDdxdQAfHBT1blc9B6nAe6wQf9ywSFeg2R
r6Bn6TPa0wsH7AYMGvR0F5h/lJNAb0cRX9BkzlA6HA8ghK4JuJrR5QBLsRERjJkp
2zBwcEeoQP/3JNcsZyShBlVrDI7XukQpzZAzfHB995Emb+HkcGIOelzpdNRqs3kQ
Yec0Bx/kwmg5mMwJI2wGZsD7wBIVSMuJVKU6uqBBnj4TglYYgS65pnAvak0L+f3L
pVTim2OZ7vhYyJnsHAl40QsEXoDmcmDN6n27TLQVVgileNLfYJ2PB9oIMmJnDJfP
ouwTHwe8d8OcNCQ6Jn67RFbOt2RKTJ2EQmwGJJ+NWKY6x7n+8FIBoq81yKkrPYno
pYkc9io0DiSr9idRynm94rxa8K2s6Y0G+V0Wow01YIIKhThok3qrSmNMPdSZmWna
2sSdT/yReCoar91ovwzstQ0L15aH7652Q01ixHYTB9prAqo3LVY07yZZi9Ulb4jg
O4/WwoipoTDoiNzCtxP/zfWndjen8fExarSs1xUmRQBDEVShG+ugc1jAMFBsbHdk
7INUzff37sPq4fhhCoNbJdmBFeBXBa/xAzvMX5iMy5+Xlu/u7/iC7NXYgTNYkyKa
vzo1cIlnqY66Ox4YJ3YhcywjNgWxc0jE6W0mlnt1YeKENsZcy6JprFbcvHTYj8YE
2KuQgFk+jS4tQwd0aBn6w+E9U4atfpVP9f8NsRWRUNKAzutGx5bdkpynz26qh0sA
ol8h9iowu4vBGtjocIFBIQ8mh4K5A/xspe8JHjvzOift9wvYXPKAe5kL2H0sjCIK
wwSivUqfzk86doI1kbLr9XBO4glyXPvEgnAm1AZzXFvZRQ8gFsmTZkUEeD37bFVK
yHNe4ny/BvMZ5NLBrVzJEpFWEbstuIVFtwoRvx2h1whi4Kz0xpyiZBgH87isQrlp
HqjfIWxp6OUroj3B/KLsp5xm67mdklcEDah7KhDlCtIbVYr/H78fDxYWcrntarFo
VJGQekUJUBi/JbM+IQ8ZqETzlTrF5OIQtFoKyrZZDJK7g1kLmez2eYtKMq3x9vCF
TWuzA4GbJr7QRI8kky2YJnmnWKp+T4yibmFKHOtmdoMG+nXqjqepu4p0qDq+v8FO
H6wEEEZF9n7iKT1sxDOV3j1m6iSbV+scvkvOicznEuR1TUKa4DfxThNcv2F9xq1I
QE+BnInbGA5HekoSlzHekci9HdwVpgfgx1eUY9hKk2W4Zlz80pFUypnIJMk7CKG2
OhR5taEOx56RUpoAB2CG2zCWBDXfw8ex9oKzFxBcvpGqo52xC58aQLpt8vn/ouYr
6Apz3UrMixVfBOcm69hO2EG3eN3q3NmziomCy1x7c8wb9nFuSL0wRTf1EkgU5RE/
XhnhZn6kGWByrcuUGRaIlnRrKjYh0u8IFEsZnqvE64HV5XIOvQFV+sPAsjRuDK4O
/EdrZDtXVwKt8JaV6BvBjOw1NFiEqbUqDyKkS1ova+Edeuu0CH7BNQzlV8x0LJRW
6pk38M+PXI4cg+qkG6BfbmwZg2dk+iLuJ6IbdOugv9SxjpnpRYX26ZKyIl5MsTHl
v7eIUFHSbd2Wb1t4ltFHrOqCOEqqZb7yEfc4kRPWOQcHiNDGS4rBGvOZV8fIbGVy
l9w59KzBVHCU0iJfankVmAa08yDluhDQBcIepWs3uVld6WcfmrXh0sroB72EywZ8
+s2lbSRPnQMZdNd18FXzzrVwVD5CbcbwoqrmHpkYCA4bZCCXAbdd51RfkIOjuzkd
mta4YL4OQTwvIuQOSr4mTcPGi4pbnTVckFoj23V3DMTrAFAfVdbQ2jhLY+ZiNQMv
b5UtuuhaVgO3yAZ6vGGPLB51DR+VDrPS2YBQsyD0fnBJTZPtajiB5BR6Ge3cMrDy
VN9sde4Md0oK1BkoIYGwIQTZSaL3YpWCDXpcj69az6U9QOTRaPzACnebBO2zafl9
eBrnjMxMpTrNaTiUzIcrGpphdiEN6dtxxuvM4Ew6YpGixSa6TqdRGDDBso8obiib
oNkFbWlWCslZ3Yt0y3spnij1ZR/fVHHl67F6NIcCa+Z5VGLuRbffjqAY0xu/te+W
SxnjdsjNsyyha4xmLCb3KSatFMRLwMLJo0O8nwOdeOjxwZnoPPfxJgMzA5/PRWSB
pYIj606uGoNkeLKiNJKk7RTM2FjVnU92osYHHBKDL5eWs4go2hSdGcH1kvWigbJ5
zALDL7208293MTcpuZKyn8/j3Cij5WknxpjWltgzpFh+cWNtVCQEvw/oI+oqTOLp
XSJ3row9jTsx9+CEUc+jejvjfvBHFXlEcDBIIuCViheGyxOlpdFtFFC0NUvRVpUU
VgdQcX2tIpX7Aj8YXIG7rJd/Vr2gmWDip28jU95hH/zhun3diply3/YqRcPYq22g
F6vQbyIgfbFv1l3O/Myg3SXpkJeu+/4cpGaVgMHwEpGwOYkarzlebgZ293r/H6Pg
TXMNINL50KKQNH5V/jrcM/3kUqZZ/o8FpqXX2ngdNSNRzsavlJ3q7Qd8Vec1AQtN
W05jj1EQKSApvUGgCW1C4VlVtIP5nRAaXEfibWQSeFUvvz4lp5Vef9JwD651QpeP
T2rBJ5YngG5Dy81WWtQdQ6lPhdSFkJCvTAonhi0uhw+OwVqTyQDRtBtQwI6RtqJo
Qc4M7cdX40Dswq6w/rIXdLxOAbqF3r/7rCyNgdj6L0nKqeCDRCJA8ICnrNIoK9qb
CUnz0PgjjCDD2pOtwSmxMj8zBUAAlgut4zzY3vr50iBLS9w3ncl+vWQu0kR/xMTt
PNw0wRRIHNY/A0yTmyQnIg0C101dM7Thc7oLp2r1/N9zfM7DOo2rc5jTwTDxbxrC
L4+VOQ/guPhzLknomFJHyqNmc7kUkMDrVdeXyeX02K4CMOejFCgWLPmrgnkC72DM
6Pzv70TtGnCo5kESC3qZIujYDWxfo4SAn1CjdxIejisYtPI3LAcCmVivL9twyzp3
5T7O0Ih2GfZDFIDXhBsGPr8OVPvppq6nQWvY/oijFtZ7gTLqha+QEdBpg+Jrlk8w
Oe6jr4rTnyLb4LV1lZTGcmYRNY1+Ug9s1LEXTG9s1stuyRMvhbk3vhxyFyOkBIwd
8hovW8cSIV7apQ1Yd7Xc3Vc8SkBWsbDN0j68+SpKuAqS6CxLBju/lwlhOt0rCVy2
gQpXEVOQ1szD7Rk+Umy/KLW4L+ISw8RFj0JU/GvWX/vUdYPaen2RdDK9qtt3quvI
loou75E11ttzTP/BFXkJhSF+jG0TNi0nweGmXccgY6MLqbhj2fZeU0n2a1QU+i5z
xu/bhKQQP1rVHau7aINLXY+ZqIUxLCQVORgVa7K5f4R5CclTFHsTuYu45i8OJ34H
yqE/giwTGaQjwqQwclueORReLhXYpsG7Q60YRxZIh3/fxxMUYrRmzhe/9ZqMuH0m
YoyqooWIDMpBSXugz/xhBvuWPQbLnJnpQuMPUgzETKhgDpMuBjCeY/QI2MtHokIG
RDL1/+jOfP/8gJsscU9AGxY4YggQXl05YTH7vxnAuR5gMyoPh0/HnDa1u3N87EfZ
nPjROrt4QBlRTJFIXmsBJtBgFfoLtKO07ipHCgbo3n0RzAObDoIJXf+B3OKUqrvA
Sg+SMsebtVDfmtYBhYXVeJE+e3/kFlRvNLLCZU6vqoOXgM5M/eRG1nGziskPbMQl
mPLZ8ifeMYJJJ0B1EQ2MlmBhsgdE3knh6+G4GYOQxBP3Ni2EygqLOXCC9fWHMfrB
5pvj+HSH8r3lMuITTsAwKzoi9xif/c5zeUqOgFNE4RC3x+2ygqHqM6koxIPc55oO
CK7PNPPRvA+2rfQ+OtG27z4TDMwWz8feANv/kpnseS8ZfvrYniFPEdicKGKaTkcm
v64y2Qka4PYfNA4UKrb+xYV/uc3CQ4UCHveyeKQyy6AzfEfc0WCYRCanCkmoTMMe
4k1iUUHdP6rHVLgpBBW+1YMYtnbF8eBh8Musli9zDIrJbY28RiC0zapfyzIjd5wM
+drtZXnPRsJ6YMgL/bexOQFfjeqf31DHJX9Txc3kcgcpY2EA2zpE5tkL/rZKEFMH
vXOZRccls6bgsxgydMICSoOYZQHI4noa/Oz3WqF6PjSEepOHydW/5kuoFA8fdHJA
L2O/oH4BSPu7lZx8g1ZKzXXam10ZYOL9NGHKa9Oi/W6LFoK6BvZQ1Bz1vUo1QhWh
1K5C5mhxWX5sVUbaY5s00Jurj+nEYAHqS/Fx87O+QrSUreFxtDt0Be2HlBdvTEm/
w1AJUq7eRsoZOnbf8O29Ii/EWUjazO0ogscZtQMflxVNINBKbPBmLfcest7mxK8T
zMD19PwO1ZURshhfsZqNp0Bsf5cISGVukTMmBLXTR3y/bnbKOAV3M/vv03iN4gmy
bW92/J4TFP+46tV4zSJlC+sxi6MrmzJ7jclPrsidLtHr61X+bJHmUUJ82fZH8d/r
tRfrlph/oVxgpwbynocIDbaqFK3/4mRLzOaq4qksnEpFBOq0KNDvSwDhZRCiJvEt
do7Dz2I0nbCZQmyzNdTiUPhQnjQfJTlTz88rEYOWKG2Rh5dYehtrxy1HzvxnyErv
qzQ8aZBzlB/PPazeEv+spCEgCLDW7Bf0FxKpoi9C0+mW8ZrPmUREkkj+VRzp7JQq
vjH0as19vd1CMgfnyqgf4zyOIxhF+C35sbIWcLL1TNz+lG+cq6oGrmsYfODpu2p3
9aRM97oIpwLxJf7I8ZGZIbm7yMKqjHMEm9FKMSnRTzdC81Zh/XLrFAsr6OJmndtI
9BJ5vzChMbBf9gqk+wts4UxfChvaL+f2I6k7N83k1p/evQhaR4gmI2pUwj5F8I+A
Vn3Uv6UMvJCPRxvx7OLSGiINLnh1nlsQgAqa4GdvGRNURxUKoSqvkZ751awQi5YK
u1fkN0cnlCcmpTYTUOlqWWVTE4uDmoR1ux3FuXANFyr7t8XSxDCsWMv7WTeQGkBA
dbXZbLk22Xusqfby6rUvuZNl4ezsjcRj8DSg8bXt96BV4wBKLdPgGlYWOseJdVB2
UX631sEP+0cEG7G0EE5DSkkRrOkBQ932r+XqUu+xvESIUgHHqLM9wuU/nm2Kg8Pu
nlRWc+ggUjBp3CM2oiBnUvZNdrycqMNr9e6zoHEieFClzBPUVW8DJUViDUyq2J+T
dipvHGq9VdG6huUqtnYiJgqxCKuIfCOYjHhc0PSIdzqe++SWd7dWT2HlX2YlAwgO
Y3OMjYNMAzf0Dikajxxq4SqCbLb0hY2Ea8iv6DE1Ily5UpyHq5f9LmziUu4uHSaL
/jGxzcYNSQh7PbfQZfkHk2nSpz3E/VnJiQAVMIYDm6wXtcCFGMrv0j2m4WP801Ne
8DsR8nWe8yD6wFGKwnsWuG3Cx8fAm/AONA9ptIA9iRzyKBCWjgA6CJodqeSua7IN
GyzzQ0E4IN1RQgBexVuzjGmY1ZFRx5zLqr/aD9Ipy1EKUAei4vJB+GRtgbCIWdH5
B7MZ/1HbXiM0zOlomyV7LNw73yBlc9PPebpPN0rPkLSyFuy4lqVh1YIQHUZJHYi5
vL9ST9CkVlOoDS3ayIYADRqi32YvhW+T37imtesKaAvPhXF4CpBH77CdYspU4QOk
6nsoeDDNi99kLBvJ0GNIj3lWX6wvAUOYEA5EXGh5VqO8oKF+/yqYbMEzODIDfKr3
lCZulcnpHeH2nuNPwSuShEesCScB/DUdXz94DtzWiqnSOvxqRyblJ8tdd5WYs36C
Ux7+AknwV1IE7enjvw6tk33eNZnFF2vJnpacq03YC8Oinw0s2iHJcV8UhUjtAqR4
sgZ1gLHWWkg1XPrMbo90IoGCqJjzpXa4UYKds+/KsyiBt1dhvNtehxAjb+6/wujV
+5hpJhGYyR4OhK3wLspIwlEykA8bkAuBughT41jiHUfqXj5VySGgWf1vqHKOB9B+
vezkKukaxgNVW/fmTVizujM3vG04DMjbRzdgNK/2EGVHvVYngHI7ZrKE0vmNIgp1
Tlw8VPI/36bUXXJL19klbGEEkV9mwxprA/I2rFRSyVoRxTF6pvjtx5rmFCDYNu6H
YgE4t94XwvmaemHE+7FRSkcR/K/MfFFd8sa+hJa4Pcm4GXanXP78vB7EFHZAJpw+
7Y5g3b9WflqWzpVGcSdJAtsPods7/AZYZguM0aLMApiU4S/+sk+PrPVmnqjU+wYs
esqAs6SCROL59iWMV3O3xnmuO+IWaJeFP5Q/cW/huYHVDksVn+TUPmn2bCx4sPcr
T8j4nC5liauh/tqRYDAxG4TVvkSrLjxG2Vmy+RZvxwcUjusISVwx+kStb341X6fB
boIu+/K3AKYs5dXg3eSaJAzKoOFmOhdO1kc0RHHPSSe8WUPkCw8WIqxwkfk4n64L
Jksieco9aYCZwMsHhnakV0m3epayFs7gBoPywlxDhcWulT4geVPwH5rw0UysFfJl
HF5N+6EbreFRrGQbb97fwAGZLJF61y6i2pzmb+D92I3RzBF7I0enPOSp0Jvc8vmh
QNILNVeWJcfQypKDRFHsRK89JWlTgPEL36Al+LgsO987BthGvsEL7tOpIcPGVrmY
8I2HFQp8/1n7qzWhL7of3bwxOOcOVc3n1+MPqw2ZR4tmjMGSK+33isqGp9/pk2Y0
a4fv9PSLpb1dMaxR6Ge+R5Bg7WfV9s1GVX1KlD08ANGr/cjd55+IeGnspxJjJOaS
hVWZgVE9hQp2cnLN94gsnk32vJkI61uIG0I8Cygd8gO1X0bsWNv/hB0VL4/JS1l5
L/MXG6yhbV9rEx7/gTNdaV64GOdw7/KGWyuTV8xexjojLN7EHVJAtxWJV+hrcz50
DE6dgmBb4xPx3K0s/1QXFCFiTt51u9OXcje03Vcac5QSaf/fHv8vkqezH3vS3Uyb
Z5s86c3gamPP4um9jAPB+6vYCB/cthU3LM9xYuuRsZ2yts3NUXLGnj00CrDFi6d8
uZzrkUplBi6nkrtahzY6ansZDEM6AQ5pk7ac8YhYbV57OH+C0qAVa3E3FMSqRutK
3p8Dq0yetHpRwJ1gBKY0OariRAdUH6TCET4E53PTvhM7FpqRrDcDDM9kQ83V45ED
icca+yBaR6cEVM7eY8VlLSVBHLLHVl3m/t2ImUj7yGRqUWt3jNj8xJsXUDRP+P63
vM0wIRRE5nCTRnR7rWEeeCj0AvuGWD3KSVkd5x6slnunugiv3z6vuaBUXlnW4Vz6
VvHBwUddq0TkfCLcJqx9gPW/zzHVBkYbqnTeTJ0CxqVNmlIihSuF78XoSeS0bAs6
7wN4EcTbXeYWrDr4b4iCCdSU5bJvzk1mnt7vFMgHmYVfSAKWGirtGMk11KDQ8AtO
U0fW6UQ6HMG6nV3VoCokiOiIjyl4hONFiTpnuU4bSoOQalzWk80j/NAG1mMq2xyY
f3n5c1032nbSb6Y3gQSPA4hiltangVNlSuAuhxCu1hNGidv3OBkawSNvvoz6BkJi
4m4m11G6FghOGjFeG3pciKGgr5LbSSEYSDN6f0ejkc44kiTgRERZCgs6StCisgNr
ktO7ARcQg1Cnyl9bpHjHPWEL8Cy+o4SzfZdjp3qtsZi4Y81tqyRn7YH0jky2OiUU
XSMSfL8GUbMYkq67+gxe6xQCYgj6T8aP2G38Mgy4F1ZUg2+jUIXLJUnFXBPMi3n8
3T8RDKwQzKr8sLctsgx9kpwgJjVm1IwJ2jZIU8KsxLcdQYpufErTmc+EDQ+kYPvU
aaRA3NzBavQGe+Wwn/Maea7aeHi2GKBuG/b0+AAntE78mdqJjgKlspXUUK5tEDRD
WqHSZiRWIMY5sSpIbjwbvrohzXhOJLP07zB3qV/6mI6/KUqin9r4aRKES1t1A5gc
XDUuXbFqZRdskyKcV/sYmQnhS30QISPjA2Nqu7g8BswTJVxdcvpuqRpLPb7YwcfL
K4B3ClprV/LMCAYDesRp6/PF7tLtsJTpT25EDBrALmaFJj58gjmjtXIWD+nxJoGk
tTmW3r4je8FnxHqonSqF8uQvwe0tftJEHNGWShP+yfMhDi3ZOu7iJwI4gnarWqM3
okW4fn+hPHsRpH4SLzfZZbo87SesZogdSU/Njbvl9srOE3k9s73bnitGc+RTFIrs
GzelR+OB1oll/1tnLuklT9AHcqeOX0s3xJECnZKd41pzJZomdWuOXM7pnA8oj/ye
HYFy2q6/W/En+tpyjRDJ4YrTrczgrFXeRTZ7c2z2yP90EOMfb10g02lwR1cxsYki
gDyVZ/GXun+BFTzjxdYJzRX9x1OC7YOQg4f+6ZoDGjI+nDP1VuM88PT9fiGvtBpY
C1eYDnZnxpJyOdxkVjkzcaABIzMUZoxjoNeiVcs8lALr/0EB3ObEYTeByT0D9haA
2FnjLvdNyLcl5rU/O0YDmFbIwT2hyKono/QEdYaYBjKAuIjIUH1HVeyvH7ZcwLfs
v++PhLmXVyP+3/LAbqsn52qbWb4QQ4GO3/yWLVSLtRaBtWBdEG7K9UIKO8mKqPc5
eCD3sFytAPrzvt+tqNqx84zDbYI/M3G77cc2IO38eCRhzNjr/7YaOeKr+n9NaGZ/
gkCHp1FKRKU1onyxP1hAjewEEJJW6iOpA/HFeuMTRUd1BWgOijOn5boCcpMGdiQi
Iv3zWzCypmgIgPX5or1DpggUcSuWe/v/UtPi2/5gEofqkwyNH+IjzBH9JiX+8GLS
hN9QUNeeAstZZcFAGSXuPn1CsP4xKJuKseYtPCddvaw15gqXbgmTD/3pMRCUwI3s
f6E9werj+LaBwvPV87IuwL2HEGKIcp2qJiW+Zgm0pMnRg33FTFiSDn5LX2QIkmfp
FgWW2miikH+m9c12eLXaXKRdmqmoRAvCsaPgSudQDyRaU5+nF7zSgSxLsbFgtENb
70l3Z3M0N+V3Lta8cEZxn0+EYv9rzgEk8LBbCZe6aVv0JA30AgiY4Sa+ClhJWJ64
DNOolAVKZ/c7o0uf+v+QHqE7nUT6/5rRP10tnNl2Twoq+p9+OK0+e2EfMIon+Lb3
dvSuo4Mk/0fwlBW2l0AGS+z2A75+i8vEMYuRzohxQ6dvSQCir4opAXjcAYS+WPle
SSi8nBEdn4BiQobT8uSLqkuZ1ePjuLe4qNitK7D43G/HkghNV7RR7bGFeW9bE5hu
ywUmDVUa/WygRXujQCAiT9qXIeI+pJcHb/gcYvjK0N9MP/fKcmbXNbYkn7ewcrJV
Q0RpbvFun9Sb/qXrHTnu4fP2Y+nrWqWP0lfKRG+YWqBqlPidBxQKK4TB9WNh+g/p
HQFDgDsr5qptmk35x9WFkpRIKXMxsD3py9Z8j7n7hQ2RtnfNNNI0adXGP4UFLYq5
rnEUL0IQyRwL14pXfUTvmZProsbRpZ4REvEiVPmr7WS5masEaDN+wVz5SuDOLIrA
vWQKXWAQ1UeEriYW+cO5o1GwaoZUXaekGnhvlxwkYIKwtTFd/l/6i/qco3S9twJv
/DF45IPyEHOvP4Bt/bWcgOno7FMCoKdXIbJULFsnLeRWF8Qb3zoQfbS42tq+2rc6
+JFWtfxsC7GGvkHz/CLL5ricnTdvCoW0cAi+Cl81/vLKEQLD0RigTWXMVs7MZa64
+9NBahQbwANuyPtX+kSDnHxCPO+5WAqa1zMSDKHLGPW3NYYyr5jDYM1nrvDxq2PA
xGnd98vRLBTflnbhmDV+Fl3Aj/+QjYgSrka1ToB0PAlKn/Gwz/geksrQWZN9gMf1
wuezeXy6ty0MBceigNj+Ncq9RRSh90c4O/UXnM4Fu/X9zZr9C+hg/9UIop5GWf5O
80RSRfd4yGYQ8nKuB83cio8cL1lqUExey5cP8Tf55Bvdy0wuuAmEzSKOHQD/RTBu
Mjp3DCWECxw5xVfnUTX3nDstlWDoix5tOSjFQcFl8PJsyoQHEJNT/XI4nflmRib7
YcIsgeh0OJiUMdKlDZGETK/ClNgIQcl6B1oW4hi6eSiHyv5Tpr+8KPKXPjoTSYkk
o8w/cS7PlRXUNThhRAVcIVMTIoWfM/pPr2NBRWw9V/BuPLgmYUc266ZAXYKqiE69
VVSXi4thIyjQKeiW5OrvwCPDoVvHMVVTCC2lUQWKyO1ewoEI+36BGPPolEzK/Xtv
t0mpU2ed75gxSEMe5TUnoGimdta8yAQGgygqMDxGYMmp8h9hAW5T4u7XxgFYYya1
Sst0Soji0QfQ/6TWyZ6EXLqugZw7X+SYXAh8lU2SLO2uVrbdVWbyGNLfU5NQUVeT
JihGjR96+AcUvcCr3crmQnHAtURTZmjgGRGtAP93+Git6ekoWahXSNrAx+659e9v
ITtDRAoaBfsbUGNJXn3fTIicW2/8vikLlRX0RLG0mQ1kODIyPfF9f+hCF4sGPkaS
7HA1HoaPYPjsCXW0+OPf+fTH//hbtuuv7qManKDVdWW3NUQyh8yDsrvIAZ6rey2H
2dtpq9XcPsjqQJJrmPi4u50Bhi4xr0m9IvciozXgwldlYuSKcA8VraNc6fOi2Hzt
EVjfaPNhN1uUXZFNoKjpuhtSMQO7q1CPC15XwPnPCrN8H/MBOlF/hoBFwXDI1rJd
9dMscxVEQYOE/78BM5KDo45SZSd5imkhXm7FS2+GSiMW16WyLppSJj4m7nki1Fhl
WqcaFDh/89rhHU95/sUKGCD+IpzoO4LrYg7K2iRhtj5mlPkWd2RifPlKCH4ZtpJ0
+xnUKzVEa8KfgkNXw2TrKNpKlGEf3py08NjZ3G/PHz5rTLEUu29Nji7WzNGv+Pdh
ZS+e/1zKvFIsIKxeLMuoxmSZnPJjjSbGBbFQMKMQnq9MqpdbNeT8NR9HTO4FcBCT
6I95mWO74Di25eHVeqfCnN+ytoufOd6wXElzlDmRiBG+KPS1/jMXvIHtYWyiz9XF
lEHWPMzyA6YxoIoa/NH2OfmcjRKZ6J38OQHAXgCHd2MdEiisRb52/ZjHgJ9bCB5G
8OG1SobgWpAmUGjL2nIHf9X4OWAWzzme/l5cOhV5GsuRup9bBgOv/SEWRyi0TjP6
EsgVs64y6Y34E1km5gajPo2nIECWyKaxcIYBXcUnttbEx0zeQeuVvBqqTEX1QLUi
YK19f2a5mlxUCvvNvsIkmzvDQ1eEaob4f1ZHbdZ3JOvaoN7ndGG1RjppC6OCmmyv
ULkHPo2koFRGxJsgnW93UZ/luUJSbDFwUvG+oATAjAMYCKgucH5Gi/CZU0vuVtHE
OKWZdiPMlvS+CO1Md4VnZ/O4oe0oDEDT2UW9cDjmn+szFRdHWrJ16bhGHuCEG/5/
y33lPELFRuo+emup3/v+5jAY0PZfM3wmGz1xKhzZmw8Aat4NWg0D1UxbP4P+kLK/
i0yMruf087mke9oa9j/1VQZ2Su9y0/WTR5MfRgNSEU6tYeKSZbG7HLwPqv1gRyog
lbtkP22GeSfajWgAsXmtDQQXWYyfz5teEMwweS4VhNrIFUyOevJh7mjz0TrS5pMl
CcAaNFTg7v4QSJ1zFhRHrs+JxEvtjQN3aPbRGic3fwYxCniT2LzoXWxyrhDb+zVS
cx0LybOKize8r3kDY7ZIgG0EHWnf7IovcxUHt+rcVm/0bYRtfrSvjQYgNR2SUu+G
3pGkiTWWKSz/95UDBeysJh6YikiZXoxIXvT1VHO083QRGDWcyoU6os2r/M41c+vW
iKPSBaYRtExg30T31Dc0b3M+XLH0vHNdhnPGOmE2T67Au8dErv0WHKovTRaVwCVJ
jtAXY/mv9fLEKg41x1bezClk4+DSLwKUFbbqOzA5vF5OxFnwFE1IMls8uOim1LgX
N0Fz8PMGBTWwfIsqtmhmh39qFFl+75Jnjd1KKOqeeC6L75vwIMn9IZXD+XIbTvdz
uHT8bzaF9GmNlxwJFDDVgEkerv4zC63hRCjPU+WQah4yzgh3o+gzCbe4N9ipRuWB
T99IYcCTITovgIml3SYpO0txUu9FxNaM6BgM2BMTG8EmhFA0R9QqoVpCiiNEvquu
mZUlqNibTEZ1ITaHzk1R9qCD9k+5yQAxWoBjfQDXZ8Xkx+bVPVZdLCBlw3TY6v8b
n4aCMR/DBCQ4kSUqCW8LXu0Ri9j05zT/63VFLbQhmgza6ZErycJPxmoNWrRrA4lF
f8oWBQUMeCCYskoSjMYLB5sZXhpaBOSe5y9f3WuMF6Awq+OW51mSx6vsogwcRsta
pIHBURmXG8NC7UB4KylgfLyw9dfqLDjY9NQxs9VMjIPis2rUtTk2j+Wh3ebMe34V
UCtp/xLzsUrltPt+vaglOwWXjctOP5fiAgjMWQD9Z+gE5UjqRt4W5FPfnI2ju6H3
KMvPTAHCg5Z0N5+/L1smbGXi+jYmDLdJmEpi5WOYr0Jr/9rS4OuYEIqZyXR0AJP2
fSRvs5oAdIOmcGob2gDcUKxEM4sOwZ2MgtS8SAqLsh2GlLq1ibHjZ59HD3Xnd/pQ
SWim/2BafVdfL8E6CoIkn3vGgPqg+aPFeX4I4a2cqf5CNg4GBH3J9jIfMegmSH62
89UwO8p/1XcsjHGp4q1Fz9a1jy1ogubXz937NG8d8jj/iFg167b4BZRD77ej4fAg
jP3Rh86ObN9F8noP7lutAzqvnA+BqFaGgr0mJ5E5WNKJPcMwdHL+pJf9vcN+wvp2
XE3bN9n2hQAORoFmugcwv1kJEIJ62s/BmTCXt+YEjkTTxwO1b1ywXlIByAZLRkgM
GkoC9R6q1BdpFFG72unu98pNfwDwbW3Fo/QbYlNOuxyUFZeCdbjCw4OM9FfNvWG6
SSSPNr73GUXX8XRYDkNHwJYOMazQUvh8vkjdVvmM+dJWmiCmy0Fkbe62URF+SiqI
nDei/rJcb7flPbDYrFpJpuADfVn7cUa5IoCOl5lGpM/9kjMW6A1YaI4llmzQ4kWL
36uotCyF6Kj/7yW7Bl4/laVWAPup0f7pm0v9C/mJH4sGaps7yxFOm6WXErtB2OEi
3+eAk9T6OZswkhRt0ua4i4mDywg39RHOzWaWPfS90oaC9dMiYmhLfWmt6sccBDYX
ar1EFmSggibB74kuIABencs1Bp+GmGUPEtS3zGhaiwZvBQFQ6cNVc4nsngd4WSp8
8FWdvVMhTq8sUi7njAEli5RHVmvIS1w1Un+C1h8A1K6yBRMaMOpJI4JvAvq+7Oyg
USCOdfNrUwbrY9dkmhGc3+oxgstWTfk+jeCCrUhEjUofLKbJD4oNTJa4ryfVuZ2c
VGmOG6CNyN32b9T6MejqzkzlZviiNCmsNkDXoQirOz7LrMC37Y4aEqzS9agEmQyf
wb4NxHLwTyrb9BUlFCuL61Ekk8GV+/EzxSXyOxvTbmMpn6b7y+gr9Alss+lvKAlS
WtEKrn47d1GAwqI/LRz9LVPJROZexww5i/Pf7gKSAbCPbTNIv8soqNanRKWfBNSU
61LT0Xe5cQE4GRIvwxy15//BaGtXJ1EJnZilcOhDxmbYhNTQMwcrQrk3oO+/TeZE
7n7JR0SGyclonvUunIjuDsCsbuHIRdJ8JAE4TOmP0G1EvxHixWG03SyGCY00Jh8u
jCyVK2M9VzY0qu5cFKTT/56pj/shLTeOT1koIzDtvz32M9NJEgye7z2i0FGSa+PK
0IEGS8G+IXjy9+af26XnZOsq0bco2rovioaOTPFtioAeiKeWxD6reH358MytWUGF
6zqT5DfVHRRpVlmFJf2YRO/Hh0OXHWr3As2QkF1vkORkqVzG9zZjanS6gkqdexMD
KX4X9yC3omnMjBirMQ8eAqMYFlk1wGLsSEV6O0CNXh3xZjbW7ZkTh1r3HqT2WgAE
l2s+mv4sTO3gsmAAQDNx+cArY9MdOcPtc3rT2f9/LI6Sw1YD1wEOIMTXJC95xiED
HbdmvwwqkWklxTLMjuZ6HvAUcrmfATqwfQl+UCT1CRY4l0J3ioulycWRlzbW3ONr
kxhHx4iSp5GIZQxDLSTG2TcTKBuC+Y93bJ78zhg+ePI8QvqFWR9VGXYFdnO+dwni
7WCTvs318ofynOxBoeuWbcYl+uBjZLB7VngPe+Ren1TVvqolbi62MUJhhrYSVh+K
HajqnvLWpFXHyttgIYHOFDxe1yGNVVAubIy1A8peSzCsCIf/blde4t9EOgPAkET+
Sr5We+tPjKo7NGokR2TbskkOywwkNY/PdRP+eN+ZLMqtb7giodWIEQt+ufKQhtTN
/4NURbKIGS5jZ9Jz12RK5GlKADUBM/CntCZu+7mr9nWptnxBqTdiFLrFhO/wnEH4
L8glG8cJ4HvUSfVyqV1f5iPgClfi8aTB6n20B9zshFuPICOJZnvXoyj8K5NZwO9L
UQk1AfkujtDXkyGljhfH4lu1LBDoEfyXR2EMowCh16jCzuy2MoKitdW7mEt2gtjf
g/L4X426h2aQrSwCPAwZtMxYmMk7GqTnWQrlvzihIO3Rn0c3NLBFfP/oBoqWLxdG
OVzdaVPegxHfIdm6J0QMYW1mp3K2HR9ReT6+DEoOxVhD05oPRAd9tEcFp1FFRD7o
I0OSjk5Z6CiQcHb031qmb2CZNa8HPsKr0fMVZ68FZIIu2a6bEHd2bO70CniNlSnT
oPAtlFIitW+26Tr8J7jPbjtlAaFfPjvOhRtYJ2CkplgD1OzPvxyI4kuplEjRmuyV
hk7bB1qPiNuVlcnkMjKdP/FRTGccI+E9yR/vJ3jMkelH/1OGszaEds+bXASrx08g
THoHl7RW5pw++y+iojcSrWRBkJQl93X4KGTksdrSBbfD3jfgiINzWtG2Kft5okv1
rSw6rWY9f8uXFgS0v/E7yP3p34uZ5RHhvj7qDr2460218PEqbTdOtX+5TE1/kzjF
C1dDzzOjSdFyTRAqnookW83oqYCAeR+SUxsYzqsyGO5qYKvPV+lBhC/Pbv/lqk/e
gTSg2UA3nLjA5iGE47EWJgmwmiEbWD9/I0EO8uuSkORofrgO/iI1mjH38CGLGmW/
ichMjFS9MFocuWHERejyUYhfZt/wLHdk9zvcsEBTFDoYCs5KfSk30wSsz+KLI4w0
7Tha3rkavOqPDUmu4zvxxUfIC7SvQJo+mQa33Yf4ZVbciHosNMscC+eYuc8XADx+
bpAaZPQfMjNy7Qn5qpoLZa/UAFQphyegJcSyfbw/Y/9h54gwr2nvK3Fm3s7Qb7zS
YtMFRFP47cJoKfn73ZsiQyFPcpNO7vZp+Hkg9LpJjMzH9yhYv6PiGMzS19RVaATc
QVDdlsg0lsmKwzU/BM+mgX2YQ/Ba4qB30wxmHY5F5NkSC/CofurOYPEVwKZRqq0a
C6w+kw6cmRImBw1l37Lhnmq6DssD51BjF7RuxCNTmQeXLGBNudyol5LY1iW9cWEP
koTNl21XYeQm8+li4ufvdmwRhEYZmQVXvLktK1P3k3fQGwTMR3nkg+VouE9YuKY+
eQCx1GOzuu43wJc4RsEtykPj3BvEa7gASnUW040qIUZDruvxCZx8FIjip9EsMmSi
jWjmP0u2BHQJw1KAGq8v0J31heK7cr4+5uHat+PFmzl4jHWbPkJRXnVw3nCWgIVt
gC8+2Rbe9y5tyIk8eHI8UkZq7renf4AWSjfW75C+Dlopyh4/m325wrhV5gz17Ads
/McupbOqPOx+AY8Xo5YbAdlxGC47ILwqOcVOhYFOP+KcpwAp3HJve1h25n8Dcecs
vQsx1RbW2MLYO50wN4Cj7UGuPKWRIvG5LzzqKaahQsXHrs4+S5mA45QN1eKiYOxX
Vr3hExlVRCywzJSb/5LKJdHOyaM+5OalJlYmWsMhi1HJSQkPOQ2+6nuTZp2ATbcH
TvxkM54jR2tr1JmV0DzmHgWFeUWe3RGfkdNq6jXzL9fWM48469gOgeVKMZ0h3uXP
tHpj1SI4e+5rFPAo3BC8zc6fjgEmgVxPV8q+Doaes7RRdlfuy8D4cCV+DuiwkQcp
PRFweFNhwV0lH4OBeW9QfpBKBgxb3bxclriG17projQQ5Wo5YuyYwTSK1t1Gkj/+
eLHG+hWKzRqx9gqgbTKVVWlAig34oHJrARNQugeG1MOtzst1tqoqCqqKXn+tdtzp
EODYhDWEqHrrKMKnIpErhj8MzhB/Kip86s1w7RqaYqxkc/dQv4VbWoyoDY8RcYLd
jEk4bTpSgkhNd8DybEHt6442KBhWEyrisV39oLIoBr3Kqfw5B6MKFW+3YTrk2WcV
T1eoorXDF9arPQvNTB4nMWVk65uF5j+YyqySmGTi3G6tESh8MSbGeM//S3K8Wr9w
rSI1golBS2K0a//VRBOw7JQdISycoorGW/WyFEx0bZCm2RwVMbLqJafEbt/U+okJ
0nEiX1sF52hQYOicKV6JIl5MgzjEieOUghcn5M5LYMrtvGv8wMx0KLPxgWQikfUS
yypEv8DMIR+Pb3PYAABLCCE/sOJmdJ4MHAi1NWuicqwuyf4qa8VME2itExSrbOMp
sR0TvvJLArYkRGaQjUPqpYlWEUbMtOvVpUhQkDwmZv7eG7y0AgxaNWjtFie4N3dL
5UO3uuk1Er0IgPszAOjyPNBMGwQi99XY9l2e2U8/8xfIZkTcK8ntFqrZEZSpMd//
/PVb4zTtg4ESTNLIHuUKOeY1caH/sU8JWo8eGCpQFpU4Ck8uy415FQfCDOHlH8Mt
Chw4cdc8qs8YvOPhyEVX39rw/m/UEdzDrjsWMZWWptK17PVYew4XLLJfWlHiiNMM
bWmlvTY9+jsy456f41+WPtHp5NF+h/uqbdSxfXp5UNcMuYzPEvzuD2wua/vCgO5F
oxAscosdoXdJsXpbOd3LhSWgQgqJDuJLij5X3cWl8J5pt7gXOrU4528siLUaOIM+
BAv3K3bq/lJQdhA/qSB8FOpcod7qsSXY1D5n3qeDEsMZ1yvKAUtoQjmlX+v4HB1K
7Nw3ngESKgF1E8jvyS44OnMfkOt+dKKVYiiY13sUyEjZL2C7OY+1ANe6phn4zuD2
8SzgMK+Rc5Bgv4+gXP3qvRiojZoqjI8GrnRGRw1g6JeWXxzHNpFqWuy5C3i9w0Ma
rNfKzc4eYdxXMgq1VV0V/YGWgvx9QofBSBr1HbE07RibCzc6yLhwedP4FYPBeB4a
c2b7AsqvGOynZZzhiZOgPpK8evtOwwKk7MdgseGVqnFNUJiGxed31ZcrLeFXG+ZH
cWZyeX2d+qD5sIR8Evp5X3eg0SU5/h5B59c0wWewXWM3AyKNsVmB8LgrTJ04g+eE
Ok8A3MHMZUfy2bc5ogZgVSzUJYxickdbq8YCKYdt259qQJ9nUsJuc8ec25Jlcmk5
/1tUlmsNHn/7j8XcS40bOemhxVtV/0wHuS94fnfnbkHXFJrCASGMwva31SXecNOc
ynBDfAiYxvlcL7ZJ7vWeLOYWtcqZmRgDiamSBHpOHG+fo+ni4IieefxF0A1uNYBZ
DeRWky4jPGkcYVc3CcAQ2utSARpfnLRD7iFrLA8cen/FM/6ziAwYHnSREqqy9cW6
MRVI3a8fEXJsmqI3qC5pqf4tmAV4LC7gLF4tXuMQni6/igydSYX8Ol5zMp8/u0Pu
76KLFcROwe0jdLfA6+Vxrbip8Q1vkHYz5sNwZNW6FHdWrrrKPjbgBanjWxw5YUC/
YVp5PvL5/8IhfxAioTwUAzjIS9gt8kPWrvnlPBpLO6y2UrM0S95zofyEI1dTUVjX
NSNhDZhV3DYhHOhWO9+HUhEDJi01CpYSfxI2Tl75cZ1A5fukdHD33E1DjmbnM611
sz8Z7V/uP/U9EQhT1pQtNLXWL3IRThmheXTm+t0zuffHbg0btVtYWJNC9RNN3fAm
YXSQq2NiyxELhiulSQh0HjpzZfyPhJ7isOj3NaU8Hs1bVS33yc8N3nnAqJJ4MOd3
891zvgp+aoFTm4sX6b1lebAM0/22ParDtvSeM5iDx+AEV4tkvaVueXz/73rPWOkK
GCAeKYDuGjsDt720p1VuOSJtwIir8SARSkyQA861UahIQU2lKm9f8+OvcjIX+UUt
ZFn+9M+Lzf1FU1/3/AwrP7q4N6uPRwd3QZ+FEb2LDztB+bofBv9IZzzsCd1aFwSP
mEiXZJdp9vBbodIw9GRfdEpmtvpHiE0Un8AkxDlKxZoKVuJ322M/TKkp4haJBg5b
Lg8iPolzrCUKJMIwrs+OqvnJgOkl6HsM0vpHI/Z6StLj6rGaj5gWJH16ThUX5CqI
x5PuR37qTdBjDlSPtOI8UddxZLed+7m5qkBbB7n8RFJXSckR1B6ikVYvr2zVCBJA
SQl35jANV0D1ObBik8eEl4JQszxRPd0jxfG7lyQP4xJnS2AJoedevefl/guMK6Rl
8H0xs5YWvITBEXBHVIYVQZSeUyH5KdWWPhhlMbYxxrPAgYyrUc40OpI4r2brUG2q
3hBKWop1gSoK9emqX7IVvbinbFLWY2XkovltW3mXDoZY5yvRRBnJCdKEbi/6plcO
vVDdYMTTPSaejZNBMQB0yxzEWBUHtzSPiD4sPFCcVgF2xSYOS0/P5QWbHF6e6SUw
fhNVzyW83UiBtXRn97ndr73+8w5ZoIm+EsaYtGOC37ibL0qKYOuzp8Lsc7X6xGTG
G0tjHaMHHzgdHzFC+uZaO0Hbc87f7JgSQVAAw1wPQUY22LRshY1rt9hOH4rQvPCE
aNAY6o3JkdjUaxAh2xDdK/S5RyQP3AlvuBd7VGVyFi3sr1v7dz4RILxq09k/glv2
irbe/7tKaPHXJ+bNprE4J+wOYMYqMQJ+1z5nK7K1Oc7VKNbQriEHSui76TuEpgd+
ZaVl1Gv0g0ilp/Gxf5s1k8KDDMpJPHsHw88TxANQjrKToT+rph3ydIr+6UG/J5mN
ZGXT0TbnM/kBuNeOH/qWIeroy+XY7MpKLThevVLy8UwF3aJ7oip4UtEJSCKM8uAv
YLODtFY/rQXplDEnre5Jld9Y0c9/Udf15lILpCc+4EiIB2G/MrYFo5HPfG5DuNdV
q94L7lTfSi3DzWJIrjV7bD4/Ey2CuTxsqU6z2e6q8H1Lb6jl8X8VKIWoHYbd0tyL
RgRghpFTW2UsXczkeMgV/YSq87BzxZLEBMYdqaCR5UJfbBKbmK/qeu5mBFji4jaU
CwuXU+Nle2LMnY5gY+/zjJdphqR/uhnrBBYTFeDATG4Yyi4MESk/+0roa9lhbPSw
63yRa6Eguno7/rUdgts5aAZeBDlRtEYAgTUprAl9J6Cy0ZCcOM/chZmvGtYnEtkH
DsqbWVOOq02jDwHI1awp7mRCIji6g9oKewbmgSmFroVIUQI9GSh9TZyPQx2JTOpX
YZD8Oss4kzj4/q7c8T+5vQMPY/FiBLOo2I/gwI10aMa+PXPpgX2R/SR2vM70xf9I
eltxZzYCSO9C1ZoGhG861W1zbSL8UVf1h9AwfAeH6Q2qrFzrm9WWw2pXk0nJEiPA
R9HheAAoL3bHB7UJgu10COw0AESkuU7e8NVkyOk4SzX4MVE8ApGBNy+TmxNXc7xB
BGAoLK4Ya8Ouvtz7tINCtxU32ieXbrudim+hXMEJYagObbBkrjaA19as0lS7D87U
9c5nVy0/Vvm16t1/PzRuFlGzsLlcefqSBFXCGyI83C6jJ0/dck+Oi/eIHRHaLBbY
8nmhbujBNWE67M8NbgVHMUJqqr/yEJC/m8aP4WZ26x6APmOG/x+FeQg9865BPAIe
r2zehjqz3Omsyp+sI4lKWtVwl3EbTRQT9ljhiTmzU/WLbb3UG4Z67K2a3o90nRZ8
43hZ5eTZcEEjpJGdCuH7r/CFrzfgPr6uCFTRw3k8ulZxzMpzVoTtLIKh7NLnDRPx
51b6kFCVAQ3xeCdNkfAufFCydL81YqsADz5Askef+xPvbcsUl6sme95WphaVWcC8
1WJVwtixXaHxZ0raJWJuEsF+5OnTI66PHgIMBDx1zLUJppbhSUZzkSuPSGl/CO8L
AtIzB7zChOdNakCu+ROQgXFel8JH6IdSMLWlZE/5Xpsoy83lciP1m4IhxHtWlSDD
jeGA5wW4Od4LnGh/C9wO+yaXkfq3tNypDcZ8YYdpvgYbaT3lvy08htU3o9wYiAR1
P8Th3FHmaM82do11MvPdjMc+ZzYEQj+vhTz9d/q6vpvYL5h0HlZmvyBfQEzRV+/I
h5+3bQ1nEA22gMcD03g/yLZqxPFIbmoBDDis+JhOTz0T0umbJfM3sU5dGoouGNLb
AjS+tUnOYqdGwz6XaMmRK/hZsRLrOlUon8PSko3pmTJIe/RPyyV+tgk2CjWiqmKI
Yi44LvLMZRNxj/5wc/TmV2lAARgDThusbNS+eTSjwlWsIaI/9STcerEx2Kik6kFJ
4EtU8Bq1gitmkv4YbA3j493PX05FXa/mzS9DUh5ZaLzjn13aq3ZbXiKkPM9hOIon
cVKwXiHKkmal0u9nj4wJikipwxab0hczO1LYgPkwSy4CN0cEIcQ1hDS8Heo12GYb
ZJSr0jEAMOMrGQh+EzkReXx2iMTviBe53AaReW75/e7rGTfJo0JxEdWy4IB+ILeu
PR55id2ahUYD1NyWH/SmG6n7/9xbamhwqqSz0gctM8Fp20JrgKSN9yYZsoZjcF7j
hibAv6IMswot+Agh4Dxzs9Q2sOwfoG6LoDkwA82GsgPx75vGUsO2nE0VT2O+QyEy
HwP/UOLtoMCLjZVBWfoP59OPhI0Qxkr/DjiJ6PbOuYbdRIQ45MvAHkAAFCw3hxsz
wP5IuV7OZCw+2GNwyiLYd3Xtb9CbT3TWwqaw6fg+QTTK0rKLqLHeQlLEdp1eUvmb
eFgRts9wBvk46hxdeUEDRMlLSTLzBQVwSuGWb66vjB2wK98QSKlHJZfaO46oHAk9
Q7XOOHG/gL0TDEv9FDoxvJ8kuDmbZVb7J8N5ELVyFrQqva1n/dq2Q0UZq9RohxQI
qkWgigHeeeUPMZNUy4oNTQb+f9fRpDpDFlhqYWF57moKQggc0jU+iNGizarRWSNv
xtVzU1v1FB40d4CiB9Z0DDYEYatas+EZfELkqZZtUTcGysx+KqVm/SFriHxvIKjR
jW4swwjRk7fvoZmg4Y0q9kSO0mvssfxutfis4cmfVD6keTdOJvS1pjme/kCST5Uj
4QnLrnxp9/7Nz7hY/+IQrJZ+6a+4VETIxzTFEDpWPlVzYWDV5kp9m+vFFwCv3CdY
He7d9fKddvmGYZDY7EWX9NHo7oLjwxVA2FaelxWVEg1N73MonlmIAyWi8E8xeO6b
1mZjQ0Rb9UWr9W++FelCzqr3Hz0WaXmZhmsvqNd0EDWgF7NtSFtmedCCKEib0Sxl
JIxw/lgh7mfWsBlXWn55mlxX/V4xH0KQNcsImA7b3vLqKgV2rUhfBtHQHk2Whev5
nKQXtq7ndHKMqDZIvvwspTQ3IB32ATEhAMCvgvVOs5tXgC+dljyVkgHbvMhCDoct
Q5txfyCyLhu1HSrPei9rmTr14kM2+3EKxvMOfsYLeyFMPZxePInjAeB+4v+77OJZ
3fq1FkFxsw28hVPtblov9A/lYQVf8/O12pXOncPtHscEr7z22YsdfD5OLuRA76t6
RvECX6RuVk1/qsC/jFkWNlFYOv1bIesr4TkDZBGMNvH0U+ue8zssdAV2QP3UnzDC
5Bbbe6vxLRBqfovrOu7SZmY5RvCJ+texiuP4CIdSfk1b1CoTfd+CtOcAh9cp8Hpw
/ni5zh5ojqIjeUBuwVBJXOS84ne7E2NsFYEjhGXbczQ2QBWd8Y4LSjEYRJPtW24k
tDKUdukDYtNPrfAfh96h2SeTjiKpxAIDSIIQyp9sHaZnsVHGauQhNI0DUN5Y1Wc3
SpBLSPkcdVvA6mY9POmPlaC+nKJIYCMtfao6tZ1315wYZhnR5lDj4xH2MWXb+cz1
OKQC6YOPKDj/9fYLW9HHJ0aFj0AOO+2dTJtYVOZt6P6wkVbcntnY2QV9C+8pmJYt
bY2qyc4iVy7P1NAPtDzLctNA8VylsP4G2ctKFJF3sXljb47rwiPN8h4tVQZbGhyd
YGj00aTR/Sy9BHClmBV6tUjUnEOc+rNGd9xC2NSsSrFb82pUdFSQ6WNbC1Dy4aU6
R8/crY4Uw2vsdl2lted/tTE5OT6ZqFU9tRQFR01I+EflmFLqWxKlOEv3SYpFXl8A
JEu4ErcqA2uv48zP6HMcDAwXNuYQEuBRHxRvkwIWXgAKgZS+JTDbGCkCOvVNLs+l
WXjNCMzf+0LaJrNXS3yCWhQm/fbJ0ymRfMGZwXfPCkCFoJ2zCpyNT3edX46o7Mnv
/It/a11ov9Dr2dM9m404XXnDtRcSv5lOgmNn+equVpx+5inIsN1ugH09iZkOg88x
Mc+ZN1h5q853YSNvdETDiA7FW8GEqTS9jGWHPmTtzB18DrJ3rlHFXOk8UkArPxp8
6FGtQFWmfqgL3VfwyPfcQ+oktg7ZMOZS5Qw7q7tYb27h0qKiNBt93w37z0pW/rXG
UpBOzblORmshPKvbNMCS79gIUYVCpQeeVnFDM6k1em0XUatbzVgFiQTXc9xELEJh
+XwadESmCeeze0/fRG20D+DCLUakkF5mEMlXFDYnrzq5rm4BaPedHbp0jJ1R5fVx
VGzsbG8Mfk9rDSH7CqfLWZP8YCzRnwzKUzY3WXbqqB5sdDIUcKYPDt69z3m0nSeO
BhjIH5n3H8Ju5WPf7Nks0xc3uul8rCT5Wx8JZ0qRpdiDWwX7fTk3drU8HO3QULjB
eidgpLofVj7JLlSXgckAHTbtrdvndAg6aIS7K+4RpXFY36pmnF2apTNl2s1MkxfL
EpaJG7M3E94b3pdRGsw8Ho+H8ZLC6K8LhWyHOBbe1gWDJsmWQU9zePr1jnOX1AUZ
lHo1m4xG5g9i8MRMJATgVgmBp8ocLSAxMZbwquYnDZfnIbo6CYpUgYWqXSb/W864
tm3aByLKf0/cRf1c0TeSWqpNohsjx8GGVkimAwe98kSpaNUd84xs53q02cI0U8SD
92HC6Hv2opc+ZaDHtmtqbyC0OwU8nQ4mpekJcCtSTjhmMmYTA9xbihnznMUkq0RM
WSgKQtbIcYRDYf49dgq1l2IndXlRNScbG6qjm9uY7i2dTkbnWptkb4j7C/WWq68K
sMhXvzoxoypL+R7EDhOYQNpqX3tKv+loAmWn7nqCbUmKocB105o8wNRKbX3hoIoz
n1e0GFDl6Oez1nAgTowoDXsYh17lXXamFiSmlNjoQ/acQ2+4e408MU9cwXEtkx5H
eTkvr3bSa6HWCximyVnbCIHa0jT37CePh715KRGCC4pRSJzAjwi0kTx7URUa5fNu
QtwMfqoQwYflpZBBO2Tmw7EVlS+8MG5cQ3fhXpCJv5P9k2jqSrRRKeqJEKMFAW12
Ny3W3ayeF6gyMhuL7qikGS9IoOOA5tVD5vwhM6PhTMsS1gOf6bISVeewCqmJTwDK
d1K6HQh8miMd1KnI/06soFo4NEei1NV4EjNyyYl4pjmKfKHwMhRgT/1Tb3C8Dpqg
41gQP4DGgZf4ID8/CcvoBgXy3ELKxBioaUudb2rOd+lQeskq5b8P51pb2ZqARad7
I6/Pymyn1Dkyo9B9NTZixk9qemAfPQ1NezQVriUTopvOY9KxPKxoVFpy/JGpK8L3
f+uAPHTht2PIJs20d+w1834Mi3MLcdnxFrBH3BUZD++Km6F2ZSMU8dmO0szPUcJg
lYs2Ic0zwovERya2ERxC1OFrKAGJVAPqqdWQNyaKXVhgJFRSVs+NRz9pcx1NKgVa
9f0gdx/4YyRUDQFmdx4FSlG58ARHIRcAf8lD6B1FK3uTGVho8eSm07NtN0CawSYt
SGj3GwjNw3XfsWNn1sT7rYS2mPBCr9HyXx0mcsVRIRK1EvrOAQ2sYnnfQOzjjXWH
lhUItJNtPkkUGclSuVZwIw9dv7jyX+D4u++hJ1nCwdiNjl0Q82Ftdq1aLbf7anDS
i39+RuBcG8E9E7jgmy3+KoFLXgygdENA2QVlRcQGiyyeNnV3kUrnysVj7dC5Ze3R
Ba4oNZ3XBvq8YJeBT8qtEXbf+p8QhhFNA9rCpm70gBtNeg4mFA/K+vrMhC/KK5Vx
AXigzUEZH20GCgUFxqm4hGdUFJMjnEvFTmsITcECItcn/O07vlbmpDkDDTgb1bt/
wcyBrWXRBavwIhmzsKrg1VQIFvxBXM7iQ8Niz+0o0BFWf+ZPCs8UcgfHJd02hEsj
bnllTLwxpClUuIzsaNdPRkf2b/FG3+ka/Ii2bdCovix+O9LKYWWVM6OjaGBzCr0Y
mcNvz1hmlcXX3AhJQ/LGp8fgcTV58QL6v31LZgeknQgM/rkbSUNz9b0f/SKB8Hig
Fkg5LvTrg0t5N8Y9X2xQrp16Et8dl8JzVPQ0B3rq9angYT4r5QcU1MVI1KJ6hNNw
dwBplnprBdfvqym9EfuICtXAxhQShQzXGqXlX0ACygJIQTUe4IoJcn+zdPAjikb2
vFvw/Up8EYlWCQmPEQPqO3JRoJPFnBWZ5xKNp3a8+JoKXwsieoBcMUTA12McBPWP
/4cDWns4HfU8YMeYktmDPdps4Gzd+K+GPI/efdDhnWiso5OTKiBGxC2xrQdCQl0h
lemdgQynuVpMIqgRzhuOjhPPAM+BJj5gNQLigC2iGFH4ZO5eW3uc1X4QKcktTwhM
ykss/+NiPVH5afFuQCmQ/TwXIucGq1Bkl0uEHbeCzH1XuMnF4tlh19V7c/FqIvqg
Eq8mgiqohKDlTvxMS1w4ak1sH+TfB1vHMbyEF84jdaxkEj7eoHWiSwC7pZJDkvlJ
q1xL41DvAU0xLn5diXL7J0yR6uaBegWH4jiHFJSdpC0lXIHlIocdFtfoYzS3g+Od
28sr7Ubn5+jlVbFZIoANO+iRY6F5LhyO3q0Apihazp5Vpsep0Shs1OyVlzg2irbW
Z8j5fLSf+ovSPcI8rUOm8j0d4meLzX6PMH/G8yMhkbQZn01Uiov/TRdtGEzlqcZa
xOcnEXl1E9nDb4ZuR0hiGZdL41rAtiFMuLcvzq0kMwchNxIOWLHcnQ3t0o4Dxppc
c8ifD3PAvGSaOIQHkcmqhGZ5yUOPpFxuVoKKAx9M2qHim9t0loKoHYdMzPajFa8A
IthaJXM2H3L/UE0x2fegb1UVCqPtKmP0UgtTgB3wdA2jxjw8zu99NI3B6lUyrPkY
p5vpFX52jH5D3VtuStGYMNRT63TqL04cyaN6ZTXXhGMObQeISEaBF+jY6NrMvFeF
5CxfTTNDszNS/SkUuKp3Zyb1rcfVfltikHrZ8KxMyHWx5h56uuwHgOQ+Vpi6KsVF
SWb1V6gpCUAriAQez4XrCoIt8lvNgONl0AIrDkaU3C1pfpPzIK3sQPzMntBi4KPo
lVqFHlU5BQ54qE+wZSSTr7p7Q9Qej1rr3tH9xcjt+uf7C9bOq5JOXS/yqRPZwWVx
UWuwDVv3+F+ArWS1davW60zuSwOSOhubci2md+mKNWq+TqV7QTAIEhLM2TPeYfHK
xAsvFwZv7zzo6uWpOH/VC33eddZAmZQ1g8vx5Ce1EUiYut2LRFf1GMFolnoK7KL0
My+XIImB9u4R7ykOaSMIIpjsQFppSWC7+21ppP/Dv7JQYl97VFJzM9zxLdYg5nwX
XbtkeTpID59+icOyfqo4SsUsw6lacxiLYa03gg23EjrIFdsy0SnNz5wPUT7YUdUK
aE/hZTVO04BJ5dkvOn1YT3TSQuSwQNryVtrJFMw34te4sK26gaDnPmhfyy1fuQ25
V6xuCbPHDkRxn+zrvclcEdkSIfArBI/0nhPtyp+F6V9j4SKqYAu6XY2pE9uQ6YlS
EoUnPdBKvm3v6V5CcdplUAE1gOXogImCgmvMs5jTKyc99GXcRK0P2UGT/p/nB6sh
aL1GqUoRGNyZGERwl3QUyyVNQwJ18GlZwBZh4tRcdtSxOGkY8pjBpLeSB5HJGWBf
VAjwLRKbyeQ1nDXdQfMvzLW73ESzmYYIomJtRc9yw06ivXYhyo6gD35X+mV7VcEp
BRhw9jHyWciy2zQIblhsy+yALEzg9F4IwNhKUQNvULkNaNUeLtBnDcglz7WUh23P
it5aRRMueK1g/TfNfb2W4VwEtQgCVDhsEvdFjnYjMrHfHxCo+5MzB0f6JH8qxbjQ
2BdlhuJznyJQHH2usXuB4ylNkuUXpxPu+V3gcdgkMdfkZveWdUV45xAV/zjGy9KI
LVMs7ch1mObDNKDg7NCxF5yYjkAq+jqze24mGWBAoLJB4yQyeus38otcV53pYarJ
TVnhXMPOn5b7oskOJrLwl0C67wA5s635j4LJ+7daJULIFULw+KjAor7Axw4Cbxi6
+MMSROGTMvouz8/OJx8P03x/xa18fXQzvU9tn8LovMCK5/VGAaaGYVkUi5T382fg
NO16uxbQkIT4IVNcVsWtxOEHoTh18VbpCJnRJydPU4n4NdSl1t03H05eoFB6ZP2W
apXblTURU2GFs5jFSEYcNruta9gFXJ5O3vAsWLQ8U7ex6xBNNIYhAAsxJnPttHc9
R/HL0V1t5cXNXMZtA5rO6fDKepBFDQTWixn2qmhBFoVI7Tt3NK0UHoalN20/Q8Vi
w5lyeFtI7TWi2ypPpEQl9rfWB8rJ3WtPB6U3LyMhlzt6vqJq9ess1AKJRRHX5fwW
9nVjvMQvbQy3SO6MtG0LxFstdqDHCXboBHe0ln+I/ZVDlwBXK083p4mE3h/R1CBv
Bfuh3ZCRZZTl9pZd4aeiu8VyTPCSS4xKsqDua5hBl2W8T9zCp2flgC/Zmfrb67gG
yvsNiiEzd8ikAwZLbQBgp3tbsvpcpaDQE2K94sWLHEVjQEN8OGAlbfHLmNCYUyvl
lLbqp0MgYXuFUNvqUyB0jOa12ARJ7rgqXLyLbtdxSkHf9ojvozwap2BhLq3yfmzo
SZGYJTESPkRtY8u5otMU5RCqqcf+p78zx2zjrcYDQprrgmyW8zj65H9SUSwN2JxB
2jk48QxVe8HcyUGMlKq/aIgOSXMdcyjL3fUp76lfaOjVvMFFZ3q3ickKWKW8GLL5
P+0dCVtt3Ca3ewNE4UTFe7JPAk9Oifn+F+7uRzhcb+2lgHT/+xGfhhDdYSBqEHLD
fWg8Ob0jNwGrAvXLIceo9gezA2otCpUAuQY0ybeM2C4/hRrxWJpQVikHq3YBc+J4
2gPCCr/YDqxKEYtbDXm1A4eTsNWzKMbfnpA/KBuRYrqV0qT6Po55LyDiFeEMABNm
lcuqwvTorfjtA2fG7a8oQV/QwLgUqd2MunWW5q4h+Lhz3C/3NViWSp5gDpeT7CiO
hrafaabRNy37zwdhZL9QS5a7b9Oi/cIWQd1L1OINo4VgMIJEDNNhmt1xONtmbIQB
95kyVnv38BoouxhhldLPiZW4s81bAtTA2MztNRH3S9MpOnOFyNAqrTtLFN4I4+HN
VLEoB96dAaYfgLIsm2zF98YSagtoEZXENpm1p3oUedhH+6WwFLFShcu2hUlo2Szu
8+hbHWxb6AP1l6l0ZOA4Fs6ZkKRXLo1teOZNeMcCvIRxHLhFMNe3a5I64UcWCMP5
Kx/sFhAxWA3VKVkmx1o5r/0XUO+fXqARES5aYr9a+Cwd8suyg+ffkrTDtTtauQLt
Ry3UeDEvvBxXGBIcWDITQlESDp6go75Q2fvWa9x4tfeMOJbCGQEjG5NKf9oQNA1I
MM5nIbUpd3nTUZJLd4lqI3ZinqXLmR9qPrNIpizDnJg6rWfCASpDdsedtybKWzkn
BLCGkUIfBiFYgK/ZBASgtM8k3cjOQOumgBKFFycD2wBasTS9rxMOqsaIG425Hu1Y
2qWJ7nlmPY+Rau74Gc8rjEfcK2tpRwQdbcWwmBbbrIkXPcRSgWMmA32mxzmGFmmn
rVjmSSaPHmV+r5Wir7y1j0jRlD3a2q7xGuqgHSKparv3aGt0Im57KUwa36iiZC+/
hrH4ENljYXj3sE2EeDueE/YAKZUtgrmcMfUctSZxHF0A3NPZlEZ3r7SIBOdT65KX
CAv8/xQa05F2Qf09Bz9dBch4WsheBF4GnQs02hpDB/eyEimGrKmqva0tEiygp3cS
dCY/iur3UT1yZJEWQiQCJhVXUWy9ektTG0NcU1SOu3urMbQpjpwaIvHHD4zmq6v+
2ack4zgjMke71UPgH5WwMfwatbD3qYmHCvsBl5J+pbNd/HBuGJHssKgvBNudnZ0S
xL4osc2wxAIZO6+8xHIhONmmAianJ6Zl3JrtOncwtdAhyAY5EF8aRzoO0Lm98sRG
Du4VzcmaW9HyU0uzJBVaDYGAUh9eksoLxgF/M6hJfVXijyAp9oVWWqHiw9P5Cfc+
h7WFY2vje3F5FIVPK4ICOcbpdgzSMlj+8+5+ZIBIjxLL2is3/UFGjHr5Z6XbXICD
JDlFl6sR71evBm7A+K5xai4ClwCFBpYi81gnWGMTpXbL3/fHjhW4+SYFInUy2suN
RgMIuTbHqFMPK7bj5gLLHTIcFFrOtTQUNLs5ZZujB/NypZ1qBMn00VOcVkwS5kRI
LbzdunSTmmoP2nGbFbYrMILsC/S0+qm2VZM0ototDCCvJAw9Ve3ch2me34VAieJ2
wEglgiIpOL01KgW1BWRcXy6sG09UALGxLVk0AvchxUoW39jBEsBrZNVhX/PIbrSJ
x4xkcFUKrhO1GJ4Wtg9ENBls9n2HiApksAmsdAoYS3XfuorWVbDNJr/w4zdzeLFf
2QdF2Y2K3G0veCqcq36DKfOrOJYRSP/r15zbhzXOmDmWHozxiiC7DIBpxDimUjfI
Tzbl0X0CV5lshhferbMjC3euMDZkqt5Zgb7dwzrPXq+rs8ME47UlvtxZoNtQLrZr
5Gc1tXBk8nUDaVUjl3/ocJ2aim7HgspdvguTUqo/m7VGSe0tVZFjCOXUS2wez+07
+xaj5ZDHFjBZ22UPO/F8EmbvJwhqbqGKlTeoxoZzhn3VF4IxNne/amDTH7N6m8iS
Ty4wn2ieK6SFOwE5Wspdv+kefOFNrJUnhExoOLbh7mYzmpjzVXdf1ctMMrQLSA8b
G0kH1X3oXAXChJgDRfa5XTI+B+SfxIXloKERcDwWCzOMawOlwJaZ+ByvHPb9ZPGl
2Cwd2BZuItdgLbv9rzNe/+H9nZZUUZ9NLOyaObbM7ieuO3FEayvGjBvMEBo24Wth
HunUaOMpKewjkPTSXs0T2IAI5/cUYX6+DxO8vy432M1uDIBQEOMlnV/BNyd60snP
JMX/UlEvqM40EkVMJp4tPEzVE5wGsYVpsmB9FxioOQ/1auqN6ip/mn2UmoqDcD3B
B0CyfwCSNt3CKMtdFiW4isixRcCYc44AhbGfpqOEXcUzeLp6tZToNvXdiOHlmx2I
S3jP1hCemOoxFy5wvq9OTAXHVX4qz8hkEZMahZEbuj8erGmmAHTkdXD3bO3IEIHe
Ip04x2q2XownpmiiKDpXWQIoFCBgpwVcExy/+pEXnTp0NyIr9obUJEkEi7WERqRj
9GDR853fEd3h0EP7cn6OyOC+rSngOJcxTQPldkgx/kkv4lDky9mojdav0kvMgdF9
hs1UuM4uhTgjuNNz/oDOQZPjWMslO1dgTGTholNaMMyOr/VDeNEOsP7ROZg4dBec
uag2TKSoe9aXanQw/UKIRcur3ZCA5EoXymduwiaYiz47+FLdUzRQhDHikdT5XitP
hoIQxDJEXo6fZrbZpVBkKEDkZAEh/RYFB1cqGKmJU9q8r3wB+lrtJ0I3FYKUB4DJ
bwuT2cpIZgUTuLAgyrCCiUCTzgrZCXt75O/7wYTb6JaB8SzaxzmC9MO8MF2QhpnU
CEIaEpkWlcZKb/4MyESJhTAS9KyU/vQzxnRv/hdoCxG4/m8JwNljYSQ6qcE5aaJX
w6uS36lXjBiyyEyWSSSeDXW6iknxIMi8H6+LCnp/xRwIPouizM+uwSxM7uVtx5aa
UQ0S334fowWvJ8BuAJHnxzINJA++EHc/aFmsrvkImLXZpm1y3uc3cHJBZDBk8FmM
Ka5evYvd2zJ607M6fEWc9IPm1Y5libvIkfSGByjViIXyklGVpZSokCMtv3jWnM1P
wPQP8MxMM6iX+G8JsUoF0Pg+370aGHBcifvq/clSqKnBFevl735Y9JCspHWEoCuX
LVorLCAX0KVT/iyF7hRgK3aaz0oHiGZDpmRjyubPHFO4NlLBHJKU94CJ7MhgdyrL
G1Cum9+j2c2rNtuPBBV3DLfPp4s22+eTvwmBGyGeIrsJhILwdRuWTEYUUxbb+k6d
1kZAhz1K+nUOC5WeP2DvlyhVibwGC7zO1xWUd5mNk+OH14bByPYz7XHFY5+9RyjB
qzGhtZtwpXDCX7BfZR6ZppggRn2hp/x/4qZ0CE6pHspjveaRMe+gGypHPBZrVU+C
2zbP5BRKPzYQqBRK4qHcKvdhjt72K888HqPkiv8l1nFqFZdyhvYP0NVEnOOM7Gpb
DhsZ6sn+GcBxt7j9aOZ/M894Uubaty1HF5zWuhIUTLHslia4fqUkMYbSH0M1aRUh
f0DudcjNPQNrVTFw7qmj9wXXnxjZ088XT5DpFlpuDhLbkEVlbMlYHXpB2m1lYIwy
MycnUt+nna//p40iOLbNX7P+fJMVftzt74L26uB+hBV5AjeYJEFsi/LXvLNkup7r
d+uzrt7KtwZAmZAueMf7UmHo+58Fe6hwOh4R3zVYE4Vkg7lUgqX5whr1pytE9iZ4
AhkRHHf3mtHW0suHvTJkX4IwgnC2pQTQeSROl60szXnznvSF+BbKaUFdTlNdrC89
FkwmnztJJEzw5VHtNnjhHvLTqgjbxiGSwORgMEepg3wuQAenPg5kXmvxIsjpfoYH
A3PRdrmc7wORzrlK5AOm9Bu6qdlRIiLwXyxUhysW+tmJ6yuyarC0gQdQPOwDDwcb
B3t9xLtS/2dGOa7bWiHYy/Tz5pnkZkPtRDGl6hhpghC/EjrxXhdY39ZLRrgdm5Kj
cDWvj1JfEA36T4bGQ00rC5TV66Iey3KQumEDdzdz8qkmU9v56TH8EQWJZKo3BlT8
Z4f9XdySP1M2vxsD0yNKh/dgBB0KZsAx9zFM2lIVPVoXy4C5HVRbMKI6eCvnCsTX
2M9+QYSuV64aGKXZFQE99Oe30B147yagJ0DxF842id6V4heKJuDbP5tyC0LZo3e/
RWTZue5ezBV1veA0EVwDjht47g6YuLloi/f8uk2/XZrr8QNOY90UEURfJ63UYS48
Tn001jEo4p2azyAqr1akhFm1mU/CpXYwK+VMWq4AD+vs/Q9ropHwOpDzk6I6bDGH
QOq7FJMB8kIz/FKNrAfBv66sweiifVaphhYZ4WXWHHYNEdgjZUGabjmfS/LM992v
egh75jBvYdClyWIIhSQVeM8FRrqSEPcL/R1LblMwFH3/PUMxc+czAQm/zbWMoi2k
Co5hG7IzJhtj/GV1ztbR6Ose5XJq44B94frq6ci6nvwxL72rAnDapymsvm1ZZ74I
ECD/GL4an/hYD5WAeZDv/AkabOc4MPFDORRgh7N9bAx/s10XF0QATyTmclWZnAHt
Yu5kLN8fbFY/WBAMuwWTj4onNZOJuVzQbColJV3FV+rqQmKqQe2opCOYmDGr/b2P
Ib41dAIDo2IjirO3bHILraUCjnY08oN/Nxtgqk1wFmW9YexN566bvHPMxqtJAAkO
mSno6Cr4QyhadSWDSBfhkuoTWxunZBJkSHTfxyacDAR6cX3MyiHyLwS/1XIiwSuL
i2WJ4wGeddLm5MhY96mTaa3If/QUG0T5/i5D36P0SoDnm0bWVJ1hdP7/cnQWuZev
YHAPtNinApidALLEbviR6Ngt8YvX4qREnzj4myrtRbumbk/OKIxlFt1qhnuvI6Jm
QcyRUi83M6w5CDtG+9YJ/eubeKQnFZxzqJeM8TG8dRo4vLPfuLbrVW2LxZkLioiM
t2C9fGL2h+5jFonfZkI3B/RHlA4GyezuDzZ/JKPw2y6PwHMb96d7DR1XMPlyIxZr
J+YCRVV5Y9A+SJdCX6IfFxj/QZmC+qEGb+wzN5D8kOjJy6LVMDbDobDqkfGR3tY4
xnpqPhmFEP7ZGvmvx58rU2Fk+Z1NI04kI8l63/i0AlD+ZgIR8XtgAOvTDNhTgcdn
F2WiwVwvVkElPOEcCw/zFkQfjctKW0S0EODMlVNNs8zMQOvnofCmuwg056IqYdnK
Zhi5JaMfPwAqy0/57y2i5ml4nQj7Ab94BGOer5P3ufQkkw8LwvkM4layjtPxuV8t
nXAkGUDjAI230Joo07FZ9vOQll7p2nXvgAiveNvk0H966hJOIvmFlJ9phS9g25pQ
OXQnBUtwm42sqnEB9iwIyOaKbmVsiW1R8xREw7UdTyf2ISkkfkn2Q4DhWCTmozzz
6P8G8gMlDiIKulTlLa+xWSKIA42YoZI0i55sK+x8pxKhHap9d1dtVfq5Iilnf+GR
t+JAfUjIZbT+eV5CAmShJ2yQ9ZSn/OiLbvkej0TwBC1I3R46BbrHuvcxx372F9ue
bYDZq28QzNxnJ969fR7z5YKcDblHnuuezRbSzr4mf0ZS+KlFCm7A8W3lO5tx4dxI
VxpZViI5Q5qX3mHhuhp9i42RedY9ulGysG5fmT7O2MDQuHZNXvCTyBOO0h8HPC+s
t67q6LsRJrAd8N5mxUUGDR2PSWeDmMB4iirSP1q2dsTOoe2fRCWxN3nfEDy5jjFw
9TxWSB4XgRdotCjZVqEwIa+YN1XgngGh5WcY3HIx+le8JQqCfEx4+HKfI1nVJT9K
c1hTsoUEMF24unGf/GsjX04/lLmJXD6A1N+1+SXhggNveLcIgsB8ZbDAgky5hN0L
9m5ZXdo2jQxSA5OZNdjzBLTo5Pdj9HPuYOZ/XjWQfXoV0RL+3UagbUCPbCDwM5Tj
aHgXWYJqqud98VLL20WAyTk0RhVzjyGC5qiVHa4Bd31pDOqWS0or1d7MOJcg65c7
dJxDTuHWOuDXgIN/fJH7T2eVDjmeP9jZg/zKhWY3FV86Fv/pr1Epc/tlhA0qjOVx
Yc7koZrZyS+ZdFwAEtdX30seGPiysV70H8GVFh7nBXxYlTrXgpuzxHx/5w8dO0yv
9Ljj5gztKk2bqSh+CU2Mah87V0I2U3IvjGrg3geBf5VJoj6pKmWuBoQ5tNFnikRZ
07liXFGsrDLzZUo1MMEE3ZfyHRClziDDCxyvQz5s1gpXp7pCYLvHtVGSNK2RDC2u
w64l2aJq3gYwLlN0PVxmMtkmVn7ALy/0bw3bzJl++HGyPqMjvqBy6JlPN87ld3cv
UC20u4V/k4yYi/3I8/FbiV1/Gxg6IYDdmuu2RJc+uSjYdSriJnunWZMMixQWEdEJ
YS0CehkD8Wq8NP/YXltOhp1Uu4XDMPXemYTojjWHWodXM51QPGdvyHSNxw1GuVRo
dQVzrmkte9VA8WANRVq76R9m+4leowq/zy/0wSNuex56z12/rWBB51ByaB2MFgpc
bHP8f5fDDCyHcCphQZ5BNCjMq2lysmKfi+IKoh1gsWWtUq3tK+JW3Sy6Y4UpUBqU
vxw5sIj0WqAh/zaH8snPKgwJ9jp+TEwMQpksn5spqS/HMPXn6vjDgxECqX96saS5
ur6yf8JPiS+EPfyTL0UCtE9IVxBFEJ06UHCsH6qx+dB2mqM+3xqBQ9To4LCwuIc2
HPpvPOT+t2uXhWHNp3p0l3whsTJ5u1qjiIKUCFCbMQaXCf8IGpPCQuIz4s2vFfQr
PpVIPJ8qmqgAfm6Xf0j3bFsp08HY5c/Ts5YUuwhgu1PCqHCoPtmrWeCLmyTzr69u
hRCG+CpNFPRijE8Vn3dqJTiNVb3docaih3Jol8P6kyk0prtQvjflgLQQaRxeDF1P
8LkJS/6UZYfLWY99K3oOP3bQddVNKAikXxI5Izp3pjUbSGT8biY/Ts7uITEPVlG7
Rr9eBkVInT+RC7qOgH5U6IRoqpAViXQuXcYxSEZa9o37ok9711RDJJe4f/3Ra8bA
5Fy9AzIS1tteHlu5JOUBSWk74IvMdjeN2ajOMg3P3cIHgp6m6LMOVMMaSbqYDA3S
jCoDBPqWkJAACua//bVWXTpcXoY4nD2NDXh4WtJ3DQc0JRgN7A/b7388gb37CzdB
BSVWyBwN8IrZoJEpX6B8oM31Cf29L3VKCgidJ1z4yxN64PG6c4zCUbdb+4+/i/WO
gJCll8HkL6nOucP+AsxWy4oiy1iOvhbU2rdSNushIU6551y2Nd6URPQoYm2NjW2p
sk94fUAnMHAarMFWunVr571kaa4PLtxTQnUr+p5x18Bm6swrCv1CefTGz7/qcrvg
u2w4hrPbpfv1oA1erQaP/tGhCAijeRiBR3Rv2DP13ntI2EGLU8Og3Zzkq6+I5bgt
/C1WTPGKFyWeUOm8gjWlr8xKb0I1rtcDIgRGzzHb6VJNvVq0FhMwLD1o5xnPoPT1
PCo5kFJn5INJpwyiHVkuW1zbSXHYIC0oymSMnnNWA4hT5BZRqqfAdGDizh95ZyuS
XFDDyLNobP1wIh6Koqxo21JGNMR+MK8DubjyVAEQWaakcIHsGbFMN2cInzyJLGAN
EIy+ii+vUa+vPU/rTtTh9zlysBzDMRDdSgZhQlOJ2fYu5LaD+v0euvtc18enOAJm
XLPJ1EL9XcV5RE9ftF/AR9JqQkpwnNOEdbzgkmUU9YIGrrslN56cJuaY8EBQe+M5
ebmRDPJnKTLqEPIVdbIHBRFokMDhtf8p6jR8J9zuBu4Qio9+XYEBjAIQ7x3hjjqv
tsjRuv6kPSQFJe0xaoJj9bTghXfBYNL94mFV/LkhtSPtumrJyxeo1UftsPUOkpdw
kRwEdY0dhUc+sdJGC92bxDjfiLLDZY3LNSBPKOt98idNh1ZAZbdo6CN0TCcbXq8p
UFOCoz/AD8x5wrYNu4GJRCfJT3mfvvKf+ssF/WZkyudfTk3y3eKoQ7Kaz+fXiCUA
xsoINSOk0piVXQuGsBRbdUhHiUwjKz+tRAteLIzMe7aWLCQo6Z7wZwZtiA9+wfUX
I5zT6wKpJdgmaS4K9R9iHhmDnSHuXNJry6pysqovNZlmP1GG0XU+e42MaJsscRwy
D3He3+JmkPFkJYJ5zSEHveeNY2818Jk7vVHaAX4DqCIOhU+eNBcgIQCFkY9lnSnk
qer5F1Jls4cbn4aK8HnnQVc0aDI+MdtNzHlQLz2cbvrdXPDKExJt2r79IBJEifYx
PZWyo4Uij3wRRKZ0Wi5nWHUYLBjjtWYKsE+ggbh4BlZOrqb3XEYy0MHf99A4MvQo
4LBiBLNEO3DTuS2JM/k+qnP9q94HWAy99GNgqBLJ1ktVNmN5ke+pV3pC+SdvAOpv
KnlJaY+2pLmdMrjMupj+m1MRyJcgrLQ0J3c8Ty8QdrgXxTYzOzGjlrxquuuK6/B4
Xif32yASD1YK2BM7lKHIlTrywhh2d4P3TpYA9Udb6qXbKuZLbLwAp1+iciHbgOJd
BEqeEqhVo32QIpXQ5ccDvodoxkkmjc+jf+mu1JeVqKhJ/gsjzpClST9hH8n+07PJ
5ifDUg0oxzl+QHFUflQhIsTLh/PpEozeK6eE3iJQyTezJmVI1gip+oI6UetMsACE
CvuXgF7mD5sDQNR7X6dbELt9pubYOl13NmO8Bcfsn4swYK/fM9II6b//B8wynlIT
lIh9RaYI57NTZEgYPVUKZK7OWHyj3R2YdTYqTBNI0AMf3rVg0LEekcT7ZyvcBibg
L9LHDVcDh9/u6qpkotqpSq0672eDzPUeGTd2dEuL6FL0JpTQ0Qp4Ob68AWYbibpF
YBpGshIf13ftMLZ9LZd0ch7cLVUSXNEiIOkgBThvhOmgDUISFudzomj/rhDEPYRJ
3Azkn23nLfT08xyXrvylMqUc8l08hIyoAMz74NPkrkQG6Gv6FauNYOAQwbAhOxtX
tdKzceEL4wClubMp4WRTOyvRpkEQcMKRKlYINUYOft8Qk0IGoOn5kLu2oYhZzzay
HLfoncUxYeBm+PIbVJXw8SHNyNGQ/18Rn+LO10qgUy7B4SJoPmuZwNYEHpohnzqs
23W7XVy5ILnaCdWWGwdplcCcTLPTg7MxIEwlCKEqlp9Hv68gM6tlgTOu89P6+4IA
ye2AbqjA1KBxQLLCeWVSRdrTtlWaf6msW6q/4cKLYsqWMdpATtE/t892MOa4v8l4
k0qr20AfQjs7llGHhG/SWxutweIdliGGGJRGiqVwt1Zmi63kFUFdE9DfUmJc47et
Y+h4L+enRnhGtCWakY/gpxvfqR1fJVvlV/g3HiIpbiB9B/ZscoLXgu68ZXuaJCz7
dtvfcbNE7NsbdiGWHFf440PG3s74H/T0XA2t5jyOnGuSEpQ3rZWscykfmz9vaA1e
H1MO2ancfjkzS3Rl0KBaVuC21PJk12pfmnx1T9fzL+4m5DdyT7kqojzXG0B0ycYx
ce4BiX/8E/quxEDJXjo0ktqE6uLt8khsTgdwlsHBagPttuFkoVRan+giHMNUh6BY
bCvyp7obXIH37dmPoKqenUxGhD40iIVTKSh8nknCeWBYMUmzgA3EUANlZKEbdWjT
zZkyVJtiioSNP/Cb65VthZ+q4TFgFOZh4QwtAesiXQPxZptbbwfIP5MqaZijdPAL
piYrpXqTb9iE2uWv0ijXoFN6E3tJxjSHudBityjL++xr99XXWoFv1Ds6cfQ37TB/
evpFXIyn1B9kKrD5ScsEscGyoUXWGaz+a3iWTI3rF5W5nW8X7fYUj5r+cMXOPB8C
P60lOsiB161Us3+uxSU5kGQeVLKF6bd2ODwwYa2t76nlL8g396EDRbYrf+PzqaFJ
2PMORYUI/TteX9NgwkNcGyi/V52zyqnUbryoYjKBh3ony9Z9yUmF/+Ark1JCBd4l
mP8/2vmHnc0nQcUvXpRLakMBy6qrhv+hUb8FDN/jfJX7E/uV7yuk6AEujOa+A1WS
kwrB89JLqCyJLMX0SZvueXi4H9JC81EZyzXpv7MTVJkcjCJtvu8qrbpdzJswoDD1
2UUBpEp3pGvEzjBJl7H/c0IPBGQsOV1bc12nWG+qD+Zynap+MfUmy1ouzqG3kpfc
q3qP6ce7M9LPHf95e9FwsYVzhG9DMQDVvOp4DRtM0mwPOJ6inCY8B7RedwZfhb1g
nw4OTc6HIfDBRP8ziCRkVnNjyg1bREwY6AFiXVd5zzVJ7PTIZlWNjscVVIJoRK8/
LzcpZLCi+9npK1cJOi1cWSUPqUCdyMLSPL7u5h1do7XPy3yVAiI3y6l2QYz1fH4M
MBFeRGaott9YH36Ko5dwBlxImWZ9YQJZqf6YQGY90iNaQ9Iji9Ln91nGZn9IxjCG
FK5clsH0581yMdDuOkKR4uQJoyutWrEAVFqfWm+JYwk3suaEQk9klOCaA/TjJvhy
PQkzdCGAxuc5E9fh+hOVC4klFHS+wpeL0YAFYo4gHNT+ZcHqb0CMQL6f4LkaOIM3
wd3+wRqznm8A5m+7GEwoo78+v7U3Hn3wdQmpOBlkeJIaoyNspP+bLFJRM9dfPWqu
/4jq5MZOKL71XaR/pq8rFwHYlgc+Vw02Q5EyYOM3iyoCebMoZls8tAqs0s8ga7qg
G54nTxOk/kii3AuwuI2ccoomCAqILC0LJSJCdcXYqxW8NCJb2WMjlvn2Gelhy75U
gVulLhJskd0BXMtrU5HoJ6jDuW4jVyUPKjxluBgs3O/vpJCeXXztHRUbFtKGG7HF
31eytHmZE/g5kscsZxjAOGcz263uSEzvUVVsuO1B9zjcsquEGf2WOSDLP4PjtyVq
TEUYfU8+Xv9rE9rUuhUTxAZSAD1sI0yTXUOMQYTB4FsUdABaoDYmGAWWA8gk0u3t
1sZvIDChFz89G2eoRCchgxbfcIBvqvVpqNJpvhrPH6SSHGCPHGf1l5eq4Ps16CHe
Eesi3rmYEgPu1EswtZKrLD3Fh8eHb9rD2W6J7LNE9Hgjis+LELg+5+EO/xo/q1i9
3gph66WFWET+pMfDaI1G2UN9H/d3VwShtbnAZgRqVDnhZ+uV9X7BOrbAc027riBM
Z90ZbETXIk88slT1C+sMqkuA9dhe9axwpIuWRajEVDUohJrfzpxL6DlZGCE/lkIp
CjP26Ul2lwW4lKLf/cwDPSWf+4ppK3waf7MOl9A6X+pihHPGmynVAKy3bUlTJiY/
T4a6avQSK8SXu3YD8y6Dy2E80CISBu0aJEP4DErx+U/j3CbvJN3mdCckRW3RO0gp
TkyzqpuhOfRPTpAuzaLNqncUBUdzEFvhMSPMGsFCFmkm8IkCD1uDb/HBHIs+DUvG
jSCNlE1We6ZoJSef5dNUDXYGVMghu1M42OTfQ+/3uhcyhIXhceROzC4wNKPP68ja
W/mmffPJax18MjyymnGro/h4JJ78iVdKbcgaRHyzSu+KUJQz/SobgzWzSxI+bImT
m3QrN3Cv6XKmRZxma3nShdhn9Vae02XVGRjTd7YGbZbcaDp/2joCvZ4aYOG1Qp+t
r7pdzPUqrQZ6PCfXwOElCdOzOXkRvghSF8jKiR1gNzngJPN3/rpOWbdu60EJ60bO
rD9AH66IjqHw8Cx9aRvq9WKSprqYxn4VU/kQHhLWjOpHifLiSBO0WDG0HU/cgGss
DT7P+n1ZmOVIACrAU8QOVBCjDYYSEsnQ0RUa0D+k4nB6ttjtskPXfOHLokowzIRX
eMur6UvODZc0uDyW+K3RfJQJBt7sNNRh0hQsZCZJd6bAXORFbf8EX749PuycmWj4
b7aj9HZQrAzgh6UaksSW/Bq6BLHWQjh02ysnTIet/HDZta8aTOGu+5vm/pP+wIxQ
I3SM3zx8wFjwkybzAnYRwiuWVT192Vsoo7R7U9gt8eNMNWtK741RurGFZVxg1evT
I0+zqxfcME3xQw70zVAmwXCkm7y6Dppt/DTApDvSF78akr2o8rGLUYynuMb0Msx0
3evWLAyJE6N7zFUzmesQ54alrT2dh4+BxndLfD7AbmFA+hXEaFS1cHM0VSkCcjMh
JsGs6G73Qr3ErR7YMzdGY/rqxNwLLiLANfl1K2sCxXROamv36cyVQ8kC1gj3os/n
eay0wnaaGqGrYpq9SWFk43GsIuNNQ2FOcuNnLP2g9cfS9bQtjtOQ5DtD5A1OA6fn
07FspKqFrou1Grji5OKRBJLofb5wUxS8bw68BCYaP1Zy1zU0UcqrT2kNKJhII34X
HPU33+SHhDufMzyhcS8AZ6OwYZga7b0N+bhalokl6RNcN+l4EP6ZFXy5O+vWZKvR
D6g0OUBI0FXX7e0rrXqGZUc0C9ufZ/8v5ElvVSSUhfjMJNKzw+5P5u/v1AfFQSkB
fj9ksB988XTLTJKa/NNnt7/sMF0A3FpeNE+VvrEiwsaSjMetP8FfKw87ERHNkX11
a8o+d9my89U+6kVcmj423aNyiXhoU6CVJd0Fn8RIkIjpiMfgmy5BCQ+PJlbjdRQJ
mQrq0RWgrb1xDa27E581b+cvvMFtCBLi+QOXqGiyehhHREmfqBxVkF57E+oF1xcq
4EQeujGfSW8/1nOZ7QKcSXArLc6w8jUD8CEEi6KW58XTJJGvwec4xgl8FEUZlyjn
fSd0QRWvDdoy7MZaJvqY/XSkTLXjyiopwBW3R3ecbo7PdBwHhQjD73V4sFAg6/bC
KsXBNr6VVXyXUjkCma2F4ZPl9kMW8VrWftl5jWA3Pm3ib+SrOqPQAkVjxQwyLpwg
5LhvtYwFuB3bgipP0e4SZ7xxD47jA7WzctLlzmS+p7UdBkH5G+tZpwR1NkNdoD3a
JlkWmbKmm/cxiB/9T/8hGYpXQ8MZPSJHTfFg2Wy8FBbAxRWyjDX5Rnk4VXJIRwhP
1GoXyvUQykPd6Y/xs+wWz0r/EFma5m7w0DIxfUgsS9d15Ula/r0Mcg8ZYVQFUbsK
FK0fqvLswMyJS40BHG+S3BEdfqMNNfzIXHxyaiBj9iCcZOXS2e/TAumoG/JjAP0M
9nZzXztqmFsPNOGUVO/9cXAiA9mnyXMxz2GlCoCIOrufttJcNUiT6SuBBdjE04L7
SljgVVzknSqdbSsSO8qMx5GSIDdplCPS4fITl5Cp3VbSD+ECP9N8ZXYk/oRvRJzT
gVto2SWz731t3z0dD3RG63TzreRAnCVVdy+QjrREfzjkYFwXCKFKOCDkuGjQy0Jz
cD1nc4jPlsSe1FnzgvVrIV1Vy0d3pWdlkTYCl9ibPNB4W0uQsLd4aEVCXh/TMKsd
IuUu0Ehm3O5vehg8NX/x4LEpI110ZbPwemipizaRWpHS2FQQQjXS2RpYjPjLOrSt
oe2KK8qwey+rjatzcC6Zp2j1qu/SzzqKJKfpsWZbiwnCpXUfDf2pXuGdkPeLR9KM
45qqqAU9HodzBs/d5Lp3GwjsE5xGubNQoe4RTlUKsogLhuz5zo+i+KXSvWEHyw9q
HWdOJTT584FbW32rQ6zdDYXFn40tmEn/nwHLysb4D7GYx0yirP4WbSvqFzQ3zf9h
Mq6LDsrs+Q427RRzdr+MYU7cQtsAft6EPr6FVkyoA7LEua1nUw1QcanTmNP0kKGd
SqgimZiGbUpAKvAx6XjCC5xBJzDiC7dlv/Ko2R9gQ9baKTFkyrYsf/R0w7TADCji
VigTexe8T+XvvP3XAJWy6Odu9oSJZoaMzo9IMqs7xsDo03q6Mm3pwYv64e7a1Bkk
DzS8Ule+IOu8K38NuBJoOkKBkkxP7ynu9SDnwDwrUMYQ40NycUVBx3Wmwx8rq5X/
msSEVgU2l2UMxpjqS/n+GoiLHS18Z2M3Zrx5lslt/1S28Icndn99uzhtosHnSdXH
vYA8+4P8Yxjq8Biq+6WEiQv1of6+3B7CiUzBp6JzIpKckqjTlqpZPqKYF33sieFy
hoP1qO1Ncmg5dKmjPKAJQz+aTyfvTewnjcYiicyo9RDzU4rOffE6kU1gPRSkzoDe
IAOdFuxfPqOrmPAB8G5fD8q/zUvcgYD+TUGCBoBV7BONOdMOpeI3NxF7aVJ5jJe0
pk+ABohXnwgREJ0rC90nWQ3dDyF2Wii/kdGRy3ozsXDRgoTU+W+aWCKjzicqhExX
VfpV0Cl+UOJICQvlxHBza4EEcK3r9z+3EKih2eucUVVXXTh0fbxG6u3gRk0drwbR
lSSkqiPehWMUqjB1X6czVPzDCyZthcTNWyAMvByc/4yuphM5gKl/ssLuRPVJ7JML
jZelP1tg4PMbro/k+lEY56rmg9avwtUQIsFnK8172gXKnEbZhOB+FWzJfD5VH9pH
yC/dSrUyJ+B3/L1NdmF8vY3KN19X1+3pLrt2p/mqMn5VYaVB3sQkDSJMv3ajdY5t
+rin0HqQKq3/kPVAlOuIt3yqS8oRHIzelWw0YW1jlDWun8bH0sJQeRA/QT1aVHw4
fQtr5Vd+U4P3XbXzqD5vubiHZ5J2ssYX3iae3eH1MpL4s93pY0mFICGPwdXPMD/o
w80QlOFnifTgWhGgx6Z44wN2L46QTzWXkGk67lGs1Kh9KMOsTeCP8wD4LhXTOcM6
e/zVUaa70YJQ3BSRHGhA6w1hQR0V3XxzTiO+ckdYX/twmgU4InQWw69b9fsL3kYn
8jmVZmJpvKcBdhTN97m1543wcqynSwn2cqI6E+sqh0LYQ1TgWVoPg+QaRrZdHUHi
gxAYhkmM3Kv5FTAvs2jcUcGBeVNqyoxVJ6uH8ARaQHmKyjXdRrUHAkXWMP0937Jg
d37hEu9BOEVmUqwVD43YddOPsfKGrFWSHCBV00i+JRaJzgmnElc2Ze6BRT0ihMTS
yFKCe6CdqnVvT05/2feeFjPeOUNnYTZh2pjCLCaUv4eig0CaWcnc28oAxQaCpW6a
TdO5yyiErcItMjw9G1BoClsE+nvJPjePXUQVxSGHVGlX/s7nKn3cgRWQJP8I93r7
CtHx7rlwbcVCujPA/7aqhQ+DqZKA4ppu2h751A1bxDcBkYpRkclMVxN4Y1Jfv9zz
GDEQKMrquecRnFNkWyMZ0x7oJ6Tm3X9K/4fZE9sT8CbfBFXgEcg23xBKeeFmz1c4
toU2RevHC6KWuL3Q7p06YGD/69GUIrnkLiEUvhhsvYKZogUSXoiShkuF2POHnJoR
FvXhSz+R2YBQYaYklpu70/2KnXjfPquTCpb5Iuybi3ZDpX6VMLc6Wfgr2i/TMrAs
bghbdXQcsvG3a4+4LEClfG2/lxCJANWh+IUNSXeXYKMOvEifv1AFaCPpDPLu6Pga
QkdgcenAAmO0BMf43SOzhmYneDkxsVvdQLoObGocZbMG0aFL1spR+XC1DDlhCQCe
UWLHooJHeVUv6bsch3SbxXS0TGz6O8inqgKfBckfQfIdmnYbC4VDlsSJRTjCobjD
GKa8uqaj7++RNNXLz1+XBej/9a5KyYidLKmcJcjORy84XumMlqXiqFtearAesgNV
rlJ4IDpWu41ayEgCaZHAYlsc4BDFTX1mDHmOQ8s8wN51OgNzyButKb+O63uhrqZZ
1MX4/ICRb+VXVqKEwIMrtqf12r9y2MRY0dSc4xYctOP4uQwdLH0UTYQrOUJ2OMqq
G2wZ7WRR4QYlzQVqfYXKx5BcS1Bku5L8801GnaiMT0DlT2l0B/7c2QCQF8zH2tEJ
LC39KcH5SIpPROgfKlk4fZXFxBIy6WA5NtE6TKASgNlm1MAPMtpsOmtZPaFLwUsW
YvZWm3AEGDJY5iiZQU+MzxeOl9kR4ykivzZZbcBaz6ugEkjoTUqZlkMlglqbC+qV
2b9E0cUgYLhg3jiwQ0TiPfk0JaB8LB/tPdIudGvLfgf8sjRKYliae6I3TFCy8G1e
n1Il+vaxmTxyIORllvRMTU+1pcqVlpoiMh23RF6uZLEkrFIXwPjL+7dlz8YfnEdg
F6N/SlqrieemmHiq7rRFONIGY67wKBbtu7vVW8832BVBHAZyuPl2omJ8LpWi6X/0
sNrku3Cc3QxbRc6ymxv+I5SZi++LPn6ZPbUrGUfnxY1uRIZA/M+39gjPCT8pAR5+
dF/1yy4bm7hjDU/NhfKI8U3/0kI9TPA9L8K8GFj5UAmhQCZa/aSYzhN+rJ39yYes
dwH+e1BMNa/kvmCnl39mpylqz/J2xT+/cSIdsP67u+VxUP16yAnz9DD+m00UaO/B
vS9tlNVkONeHPAhr7x1+1W96kc++nt95dzWFZLFCL4bkShYPSPrc8bUVYOfxjd8G
6B+y4QV7N00jum3VUbh3YZ00IADXMG7tkB84McmzyS4YYHosu5xx4sf65uFYncxJ
tnkIwR+uN+en/iuZ83wLaGJ97cFE1FEZXA58ExRJddcmGncWryM3Z/HhkNnuWu/1
YYu74+wY+AmAuLr7IK7gVPLISU8rvzsdZMIvXgQeDqQSPcpD1P2Qy2lDOz5PGexK
v6/bQxuzXMUssKdTEQKHEIs9HC2bWn21l0BowCa2Ol5sxID2gd693kuMX5enETzR
iXnJe+tZqiQ9C+HSUzvfYIpsPZDiCpYm+oCvJaPO8FKQkjclYu6uBs7avAJLgrzR
kojbvtyL/pe3f3N0X0Vxv0YOvD5cf5suJXWFN/OVINxoVLTqn8OTthDghs+GsR1N
4WOlPf3l5ySqyoY76vCwwvUPgTBZqjwi/WYdNIElFFDThsaYPMtFf9SIUX0MhJAD
oI3fD3pw45EJaj6gapr0W3nHIaBjhAk9jP9iuGvr/WkuWT15IuPTHQnHRSO+4sAk
MHxHUowK0IFKYC3v9Q0d5bQuhytqCI/SG/c/qo6Hkwwo/1Qx4/w4tZJL1g8RNZJv
74AV+lywvWXkuBcyculyM92/BnQQEQUCcAQQpHhpsiWRdzPxiYdb7kNB47w9tAcr
7SmoO9hu9sT7VQp/HtYxmdmeE63N8MZDgDltbKov1AeSlb+f1duc9dcr52QQDXHm
9dr/WvSF2lW+n8HeOVO7tiwQrecSaVUrL9VIlBKDf4D4RkKizIgxWCCS21UjfRyT
Lfyq1EtQleFf1tUiuT7hhHHutMTFskcfy7nLfwxkVQeXzoLIW+f+b6LmK2D1BsWb
66ZLTvz6h9zv+H9I8iwbxqOz93IdAeUnetRc2EXjtl1efAPC4DQRP6h84nSx8OMg
Fr0IYYAEnohCSkS7xDU0+4rWvMtPCQObBuUGsCARHfiv2c0fCAHJf1Sc4QDU0JhE
AHAbfYMLnlNxjRM5fjjrpGxE7X0E+JhoW8ChSHo2mHH6MXzF6xp74I5lnv1AqhMx
bm9koSdzPpisqH+cJ41o4ykrlRrc+KCOzD/oWBXu2lac2SQdLCDJbHjU7aGQ/nck
rW1Ih7TTHJi4OU0gHmT+kpaYtnw7k+bxK4yob9ANyMdx4IKQ+5RX5NWBGGhEQR+k
OVUlNJm+4TNm5XcDXOCk7CxNloAcmezu81HuhbGpDf1ChL36WQtcZShQLfCG95+m
VBV6rhko+aXCCU1IP8/Q5ZuAQEDX4DTP/fqu/9TBjPVF2qToRqcNE4iHC7HB0mtQ
VoMdUnpjb69csKnYLq3AtUQGT8jTcox4Uo5RteI0hli3N3J5Su3+dn0cFCCKVYTf
xKH2AFOGgssF3jtEeSzhWgDnac0pG1AamHiaPh28KXgAf+w+w9BLrNKSjLsOBMP7
hC3Kcj/4cUnluKcwbijxm7uhO7/UVwocNLlMH/28CiqwxcLLnlXAKMPifg55ZZj3
+0q0oMXYdAkYs+WDcYf/gWnkA9/XLsVuw/lP35xdBxM6CmPdfn18TMc0ugO64fhS
gDU+Rwv3NcHo8QCQ9qaxAdE+RjiwrtGaYve8EJnIe9JXsq1PaArtmllMbr+ciwlM
k2n9yCBTh03p6nkN9WJU/FPT+rObrDZ5VdNpLnNSUyadSgKBTmqj3/QY5Y7R/uTb
wn1+KC0jmB1CR7eX5nojFKpDtPhL4+geYDITyuAEqxDpIZnowXbKPiddortLCjnL
DB9YxClY+cjTnZoqcSFPmnWDrowOm0IJKTC7rGALRN+FFlYuYa6wwT32f8dY5JiL
pLFmkwmjMvMWQNPOWKjbGuFcorDIfrys0uyLmbOKM00+hjUyqh+T6OrFTa6wRGkc
NO+yPu8bMaDuE39mgA8zS8Smbe/Uby65AvXt7QwXoiAEA4u9yVvbWqnL/zdZsmR1
5glEyYNCHJHpEjZC45IZtzsyEdb78flyHpDZ3VOrEaRYKWNf1StLE2l0dDHV7KrA
6bH799gZB5XXzsommvLtxoxoLaUqsXfYSF/wykGHJ6W02Q6b5HLunYh6Q+yDxbFh
8E6Baj+m8wjRsj+Xc4zSaEQifJ+kGPmn5/TYIU7Wr+zaIi0J/tPv3cDB9cOhFP4m
yJxRKWW3/xz6VCO+NuuwRWbygkyrE5h/b0nSnjSAONTn8JUE8feCDZJY8olxd16a
x/7H4wxAUEFwHB2o8vhSwYU3saUsR8cOi9/GhlG1OZ/RXj4nHJ7miC8Hb5CPkWfb
rExev+8+ATvR0ajftCsGimHHV1wYTEaWwpnyndjmlhpUHF85ME7bxLQFjEIoR9n6
4tx7WE4bzE2UJgdEX3r8R4RexS2ALNavQTTjY1xGuDLLdLvjyq0czP4ckCKxRF0p
K5Z4b8WnbggF2kVSpzOwfJpMUwD3kNqbPctiuVY925FTxHI8yY6VG/TW7ytziKN/
wv1dFE8e9+7sQsL25KQVUqhNIqpG7St4VC3p5rL228iX0EKEBn0XpIL8mN2yhRWc
7TOwkHKY2z+/ntPIpRjkUyionwwXXwi6aqZidHub2rejlJc8OgjpYBdNbpvTXdL6
NiqSPY2VSQ5oj2KZXe6bsADr8CdD6nT3/QbBzQCbak8Lc/EXUckkGp7x7gsTXVwX
5NlyZem2MMO4qwAf7aGR7dDOdYiq/xq6aem7fq7KIrOn1ikvyGKO57WDpTEYRzUH
Ra5J2XLw+os9WbNF8fVTg5VeUAdrSCcGjo5sO2sWDYYyNBNOTAGuAo9R7do4SskW
nkipsx8FdUc0vec2L8udxCPYn0bDXTP3H/bLVGPNjwH/OXtsBugfnjbNSTY+TjkU
oUWrnn/cmQgrnJL+YXJC15YzYN23XJuslkuTcAftY84pE8HXk8CWa/uGZ0m3Scrz
DW+wOglgUcCm801WpzbpIo7fe9yZylO3G5dScH2S0eopDX2CScBKnylDMKMDB/9d
T0eTjp+gcSnMHwIZgTZXJIG0ieVyajnqpwqK9HHxB5doeOnIq15Exe3y/uf5608s
BFxaeLOBa0Zhgd7ahVWzxpoTw6w3kTzR2C5c2vHTaGowkbKGx30pVdQ5Vj8yFvFS
uyFkmJUoYws+QOCu6LoHakIJVQZa0n5hUX26lXybAk2cHu5Kp7c1kyjKVZJ66Hq3
Bt97g3ERRZFt06vOH1AVswp6o6ItdfiC207thVClraTrWokcezCtnb6sTosTyAp3
HHvpRIo0gZx/crvPayWEwZSyuf5k0hhuj4k1+9bdqvtPIoyFzm3iE6Rw3Dhiip+N
Way5Q9xO1swvxLL+b4Fcuf7bpxPG2636JAHSueLbUGcEUIFmf66qDiSq7P2zWsFc
HEC/Ycj/D/S2u6uy6sy3VUTceT2fi526tIz/11WTSGabfdotnQoAWM2DGOViaE56
V4riH0yC0zJ2A3kPRPcJW9CBd/5YQmUuo1Em1FpLkH94Q/yR09YeUJHOtWtmaGvw
bIibpi9nIvkVU/xjCc73T0dont4y+7z8HbbSU7aTLVxA1wiBpF6ll30WO+9je6tq
zUqeNGJBFj9G6qFQKna6NQL7a15lzWfVxusIwtzKl+YNJZbcvHqKVRRvjL3FoIx3
vacuJ8EZFLX3zptaCY3fQtdFv1zXpuUO8MVI8pZEOHdlgWNRFHrLHIUeLeGZ1n83
d37rJrf3DUFfehaBvnaJpZgPv4KEBwjFoPcNoZFoiNSeQQpEZ5iw+gwIPa1ammYX
XfWXNclxOmKkj58A5G1b6H3s/pO/mVqGUuDf4jZhi9F2NPoyzfJGb+IICaKoGzoO
3wZPaFo5U+hY6KwAuB4gAWVkIMyXbHlCkwMLms1owGABDeI4UE8gIxYmOKV/lznc
jjN95/W0Wy02jUydvoHAN+U6Pjnd1jcptdGauUmfsrl3JpOiD3Mk5zMzdgtM5Gwi
y7w/PTSFSzS9QmltybHr3dFa4E1P5Ihcn5zFjIykWEeDIxPApnqC88UJ1+medu2w
3bF49QI43jAFwxK2wlP6d0dLUDKl4aVJFdbs15BoSI0Yj9rJvBfev8Jdnj1mMcOC
NLqdJlqmeaDhH4oRLQchXRxF9TCEf9EURfR1tUvLIGewE+3rDkddzSgfiXBiMxAi
tutiyNC88vyUGFzu6qbIGFlfpt6vdUZuRYIvbZKMY6c0pm6EhRP5qTnXKvt3SWKO
3Zi6QmpZ5dm+ONlEXX0bDPDZHrC5jL/yBtZwUHMIm9vcV9TrKr/h/DCSFzSisaDz
UlfCNNn8zNQmxgXb3eveis4UHy29YHTQ2nuqnEzDkJK14KrRk1kYOAbji1UnhP2A
pneXzo8tnQYZ3AdZXIRWyT169ZIQfOFjzDKzMwqUd9rH3BM9yrGRyx5z66+zmN8i
11p5JJpCa4qv50H11D8xLXwyFO5r3UUsoYJafQsrZMa2WtekmvmK6HU+/kWXzzh7
Nv/pgZrzpfWYjv/NY9hdrs7zYydFZJJkvVXSo+Bg8oDKl5qBmj0XLftlw4xTwc/W
dntdMziL2ok3iupMzBcZay3PdWy3E3SfWycMg1CQrsik43xWM0xHZnXbGEhwPyMc
GsxVpcGcVCknAvM0D/9D0yq+abzelnWj0FoHRoe5SUct7hQMXHRbb9Y2476/kD04
SFdVlYt6JrtSvLVV/BknozmJ8F//0bAPt6bZLyIHuzngL9psutYkKYn2TGO+fA/F
pr61grDbxBWnIDhuUJtpLQXXqBqMo0F4W/i/6W6L1X0lgxsfWTsX+bUW0WLgssK4
PbtNbQN5eh6wiB4SMy12hgFKFJbDkT2cUzEASq6DZZErPu2o/dkHTsADr0xFnOKT
AHvK2Cj1AD3Vs7Oe6bv3kqdXZ0a7xrw16xzwqJNnJArLUSU2XjTn6u4TkOY/Fy38
XHaNKmOGVeUmO+67jzOkaeBax6uClpCefNofpZEZJeNuRLVX5nx4Kw8I5iaJNGZK
AuFsf5gIPS4aB+s3fFQwOHo2ifIQlYnGJqRXpfWhG9R4LDeopcZbsFeJ+z9EO7bA
dmf5O5kGCWL82I3LfsH5tY+zanzH1vuax4q+GlEik/IUZbFVYl+GsX1nbfxbMuos
ttXP5n0Z1ZIqi5nA9zbXcmN1HXoNMAKjK7w5xa/pRaeZ/y/8DKg48e2mltJLK48a
G8FcKBZ56HGyDcqrfGvm3AUASuElEfZrQekGAaVyE54MpF0SsfArVmR9mm9YcPlq
1wWX/Tf5xc52/Sarz5o4dLizswYk/d4i42ri+JZZglX5kcCSk9QdYQP03vvOaJqu
MVch2ABi5hAFP2BBqDhksSEWz2+LOLQtWlP+AzgZVELc8wl1sXScYwYHyueS/h7X
By4MJevEifHcniWoWHcBzH8IRI2801QQehx7o+gjihKiq3ke5QcDgeLc8UbQNk0N
IeRCxwZVsAI8rDEcbfhf/19qJhZdsoK06Gr52boH6m9kQI4ja7gW4jcRwtpLc4zQ
kp1Ul8XaAVDnbnVvzg7KwmdBGzEgo06wNUDHkOru84KiYjou+a1jyg4pCzOenD0a
uN6Q83NzKEiqHfgeTe30kB0zS1NUuT396iO5KpzB1f2Nj5xg3/z7sGli0Isv2Tjk
rCacxiuCKXVTEc/qDRp0tzsWGoYDYDK2eMA2Lrwu6CY/V7fCsAy58e8G3u6FFHa3
JBY3wVSqYS0R2mZbGw9qZtOOtA7TRrgSSfkYPZuPddkfyMWFPapO5zz58F/IIVeU
vDYl2YyY4b2OndzcqkNOKL/EA3w3WjyoPAVvjhZRmE61jAGBleF3ZyLaNG+2+PvP
cZddOvSTRrrf4oCT4OCzQTEbuqTyM8DWPspj6vcy8//1kFWHwNi8N6toIPgxqEAt
wvgraknsT4ZTf4gGnLT2V/9nhGfYbn3KzwIinALY48KvEnXmH2tABOiw9A373AeV
dIMWM8MUqx+h5UP0ojAC9DZC2GhBbi+unHcmhPk29v6sYpDtPT6SR27O7cVyUnca
ASrsPAEtWF+ct6wMZ+rP6uzy37kBK3P3hDa+Nx1wgKMxTUvo1YvNL95dQK+94tuE
mfJUjYK0krzkMZrZx9YkXfgsw119573gqukZZLR62z+M0PxKzqz8nZArIN2e5xkA
uRBHLENOmDwCXgjQ48P1sw9yj8tYsJRD2NnKhHJ2WyGc9u3nYFoUwLeKwDPxF8Ls
WHTA+dQ6g6dGB7NW8JqsbZNoi9lBroC9A6o6vYhxY4ff3/RivMMc9o2zZVJv2ny2
4e/WBFBabab6xxMBhoJXv699u8m1s9gTC0nvYfTy32v2/6/9w++vVeRh+9XCNAUL
6kswLksWplq6h/3a+q0OZ8yqmtXe3oIQtJmjcGIbmrdnkU9NYUHqZYqi2moG1Fjg
VQprcWepFR86lJVsoyfah6yW6F9QDSLati03985saV3fOF+a1QnQcxE0kFUPxd6d
AEWgTk853+zyJZ1oClStcTV5bzUHGSPcW+La+rC0elYEQaPMZ75vWK7+Z0oSakcc
kUJm4Iug+uxqLVXzm4fT93CVRrkIkZ5d7mPKJiLdbR3c3xEFOzrgdoCO5ajFT20V
eDMlyEObVWOfxUfMgl7wYYrymLF/qb2FFTBOIXj4+hwwXOMTFsMYBfV7uoVslRSm
Fmp3p3XeOcUu2m9YpV37Mj/Y4wcPfj6BWi4sUXKCQdNBqiQQl1Sry94Rx9fBLj6g
8d0a91gUWr2zvdyFquqkHJX+4mk5DMpHrgzLH7mxp/CTTsbcKzRa5XqJ7Ht2wjvb
vqaE2oxc7XlNqo2+xsi4s0eYHUgc0T05WiYUnLbx59wrRF/Oew17mlnO2H/ua0e4
5GIZDxTv41ec/SWLolVMeTLQP484KBWo9wq7axP9IuNc/G4afuAejkwKBE670wTC
SkR4IoR13gQwoVseDNJZ9/H4XrsjDqZWS+azQ5Hl0sdyW+VGHVuc10EOeXbz8B1t
LTy/IrWa5drG0h+00gnRJsDhhSa2z45qZwQ7nMOknQo6IxHD0BDzvqzXMBKHTd4w
l9KP+9LOFnLSz/fqKqfRgbNrSNkej7O5tKJwwKR5VZ6Iy6a1KAfMvrdsNH7+RSZH
RsGqTaXDVJqqZ3qSgFeuXqTh2SN/E/vS8Crn8b7+FgmfgUT6gVgDlRkn85RhzBlt
rRi+XQWXZmysVsyuW4wXVHW5gnlcO0V7Bws7ve/X4LYYFhPUil3n31ZVYl+bJCO9
7J+lj/bALmT4wlTpxGWmX4iT0+QY/ZeAZVP7zQW6CCfQIXh8fsadwfXeXS66weuo
l2QE+SO/g4sb0lUW15czXytQIfLsAvkMAXZJh6kjKZ3eL913uZEzqNv4YMMLES/7
epjl2kUq4bstlWNwklH8qUFlKFIB5/h5yunU7Ee+Du4jP1fL/yp3uRBCaXTJISe8
7DJf8UntNYv4Tiy2zHXR4zVbY9cHLsuAgpJ9wVoSZzxAukmCfPZZf7aHyK67nzSF
j/KmjFrSRe6788QhFRjVrMO/4cFdktb6Y7zG9KTzYDGpOUsaF/pB68PhGEm8v+ix
wLw1JHNsYeL8Z7E3YXJszUNAYCYHjU3mk7uzuyYyeMEPK6erfumjG8bUyydBVLpM
A//iGuZGBXCwNIP+erTUdRNXjJ53UPoDdA7wJPMUb+UsRbT1r8IkDI6oMWQixP5Y
bjNS7QV8N9vityOkULC1+5dOiYXC0aHIPz/KGOqXBxWdxoH5g8tNF2uFk0n56eiv
i5+vQVteEPtw8bhGbSbOih8IoZCC6a9EuP4aOSTx+tgnu/wxAvdXx6qaouh+l78H
CnTq/iVE3+NTQO5vDK610ynDiy4kOeycnxk36BoIKiPVnlmuOhRn0byu5bMSsjpk
ODnpVZ2gUwn8534t+Ae1ilBDSZ2K7JdNGXRVkE774LImlSutxvh8cQqBvWr3JGEW
tQ94F0GQgd7IKkWEmuI/rLza6C61K187+X65QjiPpgsvldG8jeR7id9mcJGbbIFj
EONvV1HZXN+0N5kIDy2zZrx3Jga6/TO92ax11bse95kwcMg3nSiXmruwnwStfLPA
ZxFFzDOBUTsVeL6XANbUXOYvZv5+WCHmbkT2DPHash2k6FVE6O73Lr3zoaOfU25w
WbsZOAET72m6SnLQ6LiNaUQrMWx9AWL3LWgpjESIXSFxoqziVRgVhuPkFUipoZJh
aKb0ixc5Om7LGtNriLAZnfwwX+obSCRVwXtZYEmQu/DyEFF5FF0HM1kfWmm8E2Nu
N9As+cY+lIwBalD6HDhOCW8exfQpjeWnqt8M23x9pPkE3aXRTK/KJOy1bkeEghcq
cx6i2BN71kQxKrJvMesxVHLgx6nD+dH8y4Q9zATBJr3Sol7N2CzZ+WNWw7YALaUn
FhrZDcsr3f9sYo8vdL/3AeuNhtZNxxiluCZjLQNJAaKkTZPFQpLzBy7mMthUs9IM
JX3Q9p8iql7G3GIJs/95FUTVaWBBF33eSs1l2a3YuT10o42cQfN/wq3WcYVndjQW
1p+7XCEzgzDKd0VxaLntPqVDUFK/pKD3pMc0TaOVLRhgvYWnTsRVgzcYP8bbMf7q
cujfpiIWjh+6uDlUmzuRQyxetbdc9HNOXlKKbiWtHUIu5cI9nP8XSv4RhLQ6rEyq
njTkYb3LdPHHMLIYNY1FEjwtE2ML5SDwJ38Ids3+xmJNi+g+uMYH6SujFE76LJBg
pYr2oEKzX7GtU3T1Lj1VrBFOUpCdx6OtzvC+/BZ7JuNUa+ZUklrQTKmrbP2Xzrx3
h+gpCTYmntH4evhlLiik7k30Xaglvx3m2JowOOg1XNLJNHwXT1RvXehEhtSjsnTZ
OJEQVQOVitlrg+CVENK3oEn9/cwX3qlJ9yJ1NQ+VbDcpGpy1aiNlNe7Nam0sL4Qp
/NuLqriTRatpglc31DDm2efSw9lLxlT0sWuziZNm9vdMwE8sUKsLn/u44AEAarcw
N3Y/CC3jUcl3UyTm2OR5g0Je2dq3l8rsbB6uv/FSU31tvhHMVZypuNF84HMD7BiZ
QJaItTWncN9K+B39dVrjwa5C9X4/yWRpY2hBdMwhcIJO49tXCPU2ZjKG9P60Y1V8
izuvS3vVCHSmA8v1qVbGuNC2du2h6hgjA93xT6idGVnXWHoVB9NioUAZrxJkj4Rc
8+BEYqJDA1bW8HWXiFM1WgytHbysGVf4b0X10HU13boIPmwyYa9NwXG1NMvLVzHv
VKMEHxuPEeR0lmlyXTw22t/5F2vBl7QBPvufiHNbMR6Fs9AFnCm8vbUF2Ubtasjh
1/kIGf1WIoZsqyHKWjGa/KV/emuCoAfOf7vqTK5jAEB1UMoMUEf8eHZWpUFoQCW7
yYHhIyHC2z6vPAgvDzPEoE9IPD+vMfCvtus+qA/ecGzYRwnl6iQCj/3kZbRsqW4s
fccIk1hqdH9dEPy/LvMOJPTyolplKo2QJfSANk0jGZ1v6xqnx+Hh1VMAkJCSCqBX
k6k3CRDLBealXtWNmOC18EpMtpt0Ozv1eySj+pwVJVxpjQlSHi9ueito/rV+TTmP
NnmwJPQH9EJFt/7tIcPjUK8G7zFxO3rPF/W0/8U7YWbzXiUDU9ZSyaAdqqitzLnI
2NjGDhtzBJ6+gfFSYCSUhKDN9YymbRcpnbIKV9/jJGJ569SNJfqPjBHt9tda3t6x
TZgWdd2UKelz8Vmj+4pjwe9TheZWdHdFeT7rDNTb5/s+/9DDQbay7sJFmnqrkAa7
LDSA65wCP7sIdlVOukvUxAkSUC2zM8151Q85+3iE6NfUn/Dcw+GbpZVL+nryG4Z0
6Vc6skIJ2/qPuwmkMYjUpyVEBYis88DziQhkG3WpIJ0AKttR9FYzO/JU/sIq8NKP
Q9Ey6kkKvYC0Y9tBRBPT/lfaq1bcRD8juJ7SsKktcKTLvpp11HytEo8yVJXEX8iS
sWfXLspj/5CPig66papwUbAx11Z1jisSocfESAS9n1Shc6LmQImtczVK1wm69zJW
+9gtWs5bwCuo7WhNQgMAHdeefV//UpgIBZ3KM+/XWGUHPAzBjgfdvS6+yNNjtedt
6MVmKvzUm+My7gbgvjQVAjJ/4W8FwnvZ/Bvs3b6/3ktgG6mJJr5R2f5/H/QLdjBr
FfbiQ9yFjE+HXrr5+NVINRl7QjGvKRIgZRRO5DPllRQyqPLeikGOiQ/nq1J+2qwc
+qEHuEWDjGZ5cs/vTvZ73h0MUqIJMGNM0mcJWdKLZmzX/BMlGuKdn4MzxRhXUAR/
Pfg7h+1boQ5jAR9PpzTmdHpWsjZM2C6lubTVRBjoWQ0CyQ0iRMQmT6kI2XNXSjfr
0o6hVn470agRSLMOjCcihhHSqX1ynKX7905Q35J3IiePGN4kezYpyNt1jjHsd276
YcC4GhylDGpkIcSqO3TE7f3MECOQsgyqD9FB2Kfju4Xpkou6/5e3Vp6nQbfMlbyR
UWO+RIo4KjG0oBBY4TTOuPsa75yayATSIrKjPpBpa5K4/c5aFvU5YovyOnARKu0s
Fe4ffn6u0CAR4VDj1/yrwvG+FuKxSKORLOJ70yxn4PgHGNhVj9odPdqoE0FXGId+
Q/z5+gYkZaVTiQS+C3g6pUjagPEsZh3jPloeniu6uOb/4cGbMmIrIrwStbtauyEP
vivvkkEGDw8q4gC18IDiq6kLwlWDQzbnsmdest0pPw6v6D85TY+nLI8vqc+OynCl
A84xqUfd0KfNr6XMocHo96lO++KtEBARooVh/kYy5wkJyNj6T3oY8EsdUViziSqD
+nnwr1QmA/9fZva4M6NlMFABii3huZRxotak2RsAh/lNP8dF8nfMvezV02CEEHL6
anBSKCPGSqfITRvE5R+tCA0ep85xRMW3eVHU7kOfecxzxOFZEyuiiOHj3Va2UMum
oDfurCAtM8+PONglUEYo2vHtAdVsWBWTv8jNZsoWUyllmuSuJRAbnCsCao6ByZEn
1wnpLVl3rfE7qyeHyr5TGTtjzgaVos/7j1GZcXGWTh7BImcFblkqWekdQedtDEv8
yr+VzLEeqYFlt3qBvq6v1qGXhtNnmbvnJnVp9qlvZcl1TrUunQHPJ7wk53G3Obig
ZyvrbMFtwYWNOSHuAChyeGM6d3XynHZkk1Jfeol5q2MeeKMYu7y0zJCXftsTzR1t
8f3EzXY7LWKOMi6HW2J9U6tSNbYOxyShTxTjz1HJQW5ZWVCmWD+A00xfw0mmgeNH
KUK+1eugZ0L18Tw0MKNq0bAMe8erOJHau1bpvMMEedX1Geh8u5kFpIdPtXXaDhP7
+wj9YqZxyT2Els7JnTHzH/4ADkdXAK75x3QB9qq4qTPoog456guqqcBmOAiAt9lM
rWvWsAl47JK1jL8RS8fZSvUHMzlIilMLGSZzbOABI1iLbavzNfUrf6S5uwSgn4nG
76nI9+lF21w86VnFZM6s7oLP4YjHz7vPPIVfE8DE5Vq2UuS56iH9oSNI/fFJUbA8
ewu4c/7i1SSJgjIrz+naEYFr+JY5FSSatcTzu9C3wTMSUSwONzsKszDW726nUS/r
Ipthd4jpvxTxfdfuCIfDyYi+jG8cZRpSd7FbwD3udtZsleO1+4IfuOWUJDSOgAoB
LpTimlz9QItmjxNrU7VNk6If+hoURjiPrUc8Ps0JDkiVYTcJp8OfHUH4K+qX7usP
NGIiQyctwuAVzEj4U/mxzHMqcJWKjKb/HRenj/Y5YDjkIscqN3Aw6DsHBUv5iRks
okjS63exgDYZ30eujL4yjbBp4rXoJY9z97qHomhXkaTz/RJp+gkmNVlw90UBZw0M
cOFSOJj0m+Awhm/+wLP6lCgj3XG3nzM4kpEyL8utD3mPrh9+2qUOSp5edfhP1af5
OsdEE7D6lpPg8FvtQXu5hUELHaVY4FWHG6JsUwku7uWOcbVMeeiF7MSjBt+C1UQh
q5fShTD/3yIsl1EJsAVGF4XtyQwZftR6mzj9LB3XUXJeYwBwHQUbeKsz05CWLVQF
Quy/3cowOIGJgaYVebl5vOxjD/Vsn659CWG61xCc/kuZUjTtEtJlW7q4CRiYlxtG
dUQDVk6MU4Ot68FCLsoRfzd18CP2peAFT+0wXlWPdEh5o55NIRg15uJkckMwwdoP
6RWwK7+T8DpfSuNwUHtVFTMe6T0blx8IFtfAxWBaGWh/H3Xjntic54o3W8r2eg3A
VOPdwbAms3kjeVKsmvWUqz3u9+/AhrrWeOwsQdU3WLlqyhVqPLdZHzpi/koJ9WIz
FcETSAy+LnnNLzxtz8wwKG4abPeZGFKMLtPQBxXAee38NzfRt1QbzrDYGWH2RQGD
zvKO+GjmThM4WAe4wYUKbI5ZXua+aelz4T1kCWGO32NAgKx4rSjXuGCyxwD1gabg
ODbm8gmYwSwsOhybzdh8QlyUFHD4Hs297NUERPrZlg5lOJthBJskCl//wg8BFpWs
/THuMxbt+eBmioy1pvIVQQb9pNERAHqsrkdXqYEDiSkCkyWCvdNEgUNF732ekEAi
YdL6Q3ZF4F9nzpU9eD0iKLW0eOqFeR7w3mBqKNp6oWqy6wF8qhIt4IupiTqrwxmC
b5ZDM227TW1TBqIh73ulGiAIVMQqZgcP86Gn0r6dnBQctbMtTKVAQ1HFxbgejSWK
heZjVgKIrrytMjJokWhuDddym8TjjMYPYsFBorhXdHTLOyV4ZvwNOE4uEWsTKI0Q
Z9F1k8nQGnUw3L5t9ockckQQ+4Z24gvTmgb0OymvCLtkk8o+MzGn0QJI2CuZmFFw
J+0nyR61/31mhf6/rHjrOzIpJGxp4uOUUvRmtKHgrdpPSNQL9ErHXvTw3MtxYMuh
z5qBFjl92ZZSCaLCOlgjhAUbasbLYuReoNUFWuua/h8rp6p7nnRjDCTKCNuHFaJk
uibbrwPeNnv9bSH3oGkGp1w3TjJN6PR0fslJtbf3MB8G6WoIJsCytxALPriQQqsr
WNZZIOCGrf4y5Q2VIIlG4ieWdX4qSG4DsDsfogEhM9KPYwvlWjaVWzU0e4cwKaPP
ilQq21pNUk0Nnb6w2Ta1PBw2jaTR8rzKXcqd4GBkRvreazZUn1rXZE6leYgYux9L
GLWuI/pJxm09M6y7UqbPq+K90MLjIIokZLvjPNBoJvHWS26LSxJwb880cAulI3PH
zIPBowrF1zRltCTj1qWxaq0XGM18Px/vTBGb0/8YAflNeYY/L/lsENpWJw8Hd73k
kZp1V/0e4U+2LTfMPH+4KmE1PRCJqAxM0FdDK32fPULlM84v/Nzvamtbg6RIbl7n
TFdJHbiO6ZyAz/yoh+qt08XAal4uajU9n17AEmZ280YHRi+D3YhonwUV1j4CRdsm
O3btbh5fNqFF02zFQGEyBG/PIkupuQQeO9t3jAsS2V6O1qMg6qkJK9ww3qK4Iufb
JNpq0l0yNKELlJ57WAtlTzCqOqlX++OUbvFG9yrcf1j3CqwD2zI1Cw2qMY79BZsH
e4VKDHowFc493kWCgZYRxCeG3gTV0+TkO8Hug0JqITabD6lr/0Q1yQ0DaF8FGEc5
2NLT8fdytl9Nr1hStpE3sj/0awSUSVOOfhPdPeBsMfb5IpX+jG6BLv/qOFtatLLK
XSgWbAg2pqp8xCeEFT2FKle5c9HKCfggnfAcpltxWJiyuNZk4/OSU+t4rpf99q9X
YMdd3Yp7H+qUCE68L84CvNq/KBQiamaGn/Y2uFrUyrisrO4QGbEsBzKipyM5DN52
AzS4qSxDebxExxYQle3Cp4Fk63T013BKutLLNbkA/7+H4hYKcQSnKsw7dGFlNWn+
wXL6xPKADmpliXh9VuNo9c8EupCojqa0kz/3jasuJzv0hV1f+4335wbUa9u1QWrL
NasoZ7fpL98OQSXNyxwc4Fk1Cu1kaQlwOUIkgV3mVPm4JHul2u8kvhmOhmISOfXx
9l9AzhdQcgG6Vw9uMTUAWlyfatEha8iV8UB9yXqbm74gGO+VMozm2ZFY/UyGCJ+C
uein0hkADHzWEjvn8Jw4zHuLZZUgPMoBFuscyUSmPbqqqc2NMz7r+6CJjUiUUWl4
yNjg+H6SU6AjYsvTOtZi6DUckBTxG/bWw2jGIfBWfTt4L0m/2wV9Stzu1XDT48qz
+kHl08HM2sWP20TL1FitzTkqru6ArbLv5R4wakLUqJY2rs7KLR4cEhvNBlG7I/Gw
s/gSY92AzJBc7Az9baILjw9pPehpZ637xeL5fwcOD2JEiRjSmukCZRU0L96C4qzm
xxzhAHG8QcX4fC4Q0hTSJgt381p1K4Lk6JZ7z5/QyzrIi98+Y/SLhh6gHw5utwP+
SrswcwomynaiptzZ95atABqHSkfq2Cex3wd71lD6Txubfi1c0kAfIh1GUDcpfoh5
enEzPeANNnVgYxXonar0m+CrkkertPKd+A0LY8N1zrDGi72q7swVqNWYAFuKkwrq
CJ9ukw0Es936PMS3f+3vuxyWfe4bpPHgJs1VOB85bLDCx1A73/0smraKgIj3yKke
6G9xijXkOUUVVnd9CmUGtvkwQZSv3vyKOP4dr8Z7bHd4BbOAQkbLpg8yTZc8n0UK
STGkUVKFQDU93uCWwzutK5bhc9X2VK3X2ZE40xcDwCT0DL5ps3AUVrVD+77ulaa4
x/MdFsrkbKkHtIk7rGXE+Lu4RQLMZbmZ3rpcBqqwQfSUFODy7MVBFwg/MFvLGmM5
tVUn1Tx3iFawTLL5mFIO4Aj+Er6WB0B0uXQLAyhHpLuePQlORWqcKImGWBi4C0jb
ZfXsnEAjNCPc1dVd07rS+x5TXJuzGGme0HqhSce5nvMguyjGaT00e94bCo12AVFq
0R7GohJ1MQmZjzY2PvvyEruj7V4kzFP6rkO9ZVn6+gNsL6iJPWRBgcSgYaQVeS1g
MT0sfox4oQsRxkt5jEF/hJaYb6B5XDhN45AW8Z75KqGMzqFV1i9ASfAZTtYo28+I
Gw/DbdpIhYBwOaSp/GPWKysuPb5mHu25u6IZvScCAibzK4EdQpr6WfarnC7VMgye
NhTKsO6YTBoNOiwlmmE9XvyMGzaT+HH9oVDhqTKVT4LTVuSM5lYbwdWtfWIl0za+
Fnum/P+8A9PpRddFtY8c9PQ1+fdf5vWEvrPAY94G+5e+B1xur58B7xVOOTOGy0fG
QIlL1t3bk97YdJfM38/pHjwp0wWnpzWqBZfDHnINEyyxFOJdcoznbt+St7v9bHqH
65JtWGV+Lnfo3HldpLeQcQAxLNQ06KS0uyvpgglu408xRch22n20I9g8tHBaEj/E
CmvE9gUeynQUIdYgngCbrKnodhPk25nX+hRs5dCjQNNpBZvaokJIIv7p8tqKpn/i
99NL6BCqY9LqcGp1p7fpH/dWoA9ktQMKwSOXmFZsC0wq2yBvoBisvOqoAvhkOvMB
JInK8xdBW4XRspCMPn86ynOC4cnk9HG7XiDqUk961rEHBLQUpA+HgUUCTBYjYSwj
+5D93D+7z2AOYFJ868pl5kQ4PD2toOk+05j4gghx6WZwgmu/PM6agKiZpmbcEeUf
0GKU6LrrCGCrslJzcKiKJkEutEWXS3o8yhWuuWygPIyed0TWPR4me2Qra2pCd8FA
mNvmeD/E3RdYcErWxRpXD03uvC9TqMOfrIzbMETf1jXHV4kjL7WNxhEw3zzZhu9o
FNsQZd3qs5NLslaF+4Jr9J0fvsBuMVKLFJv03IAexg3d9g/osSdSJxIYjrZ3g3x5
38/jU3IlGwHOVax+w5iD1O+BUID85KpTdxtHI64SVy1sNxbzqJGJXkPNZ4SqoP3f
N3hjQM0TtiWo59VIhqJx9SJI+xpqh6nxXeRImGcH7NkqUGY2PyLbwCzXRHwQOMkp
iPlzeDViV4S+0OfyJl7z+wYEaV6tvnhENY0Y8/FMbUsUcRPAprq7jsZwP1RjPSBe
zO4JsETNbF1GEcGynNrj4FomT/mbbZ5iBVHzCMIqcR8seF3nJ9EmgB0HrOzFJV2e
AlHYN5Q7HxZ1ZJ8JRec3+eztOjBqhyWbh5fG9vVzW5Ck0xJB3AH6T2Np2ONEHj59
4n9NNYKi/ilccXBYVQ/i5O4wV+D90wqieroHu8+JTpcjTJa2bRnOW19eJy27FCCe
FrDbD+FGoJFISorj/SLTwjICTVNhiK++mfzfv8CtsL/661dgwhIjQKOmZOmtmpkU
sv52gv48oPOVMnHrsWISMwkH9QhdKAeUWC5Q4HEANyVaD19P1gMoKHZ8ZfKkL9FS
ewxAZW6V7Gi/cNJK0GB3IxD3L6v5HL6Q/m4Nfkx7xqQ0stF/esO7o8Nd9DFJ8R7r
arhPdgzXTnpPrXTLFlWRDnP6dxr36cDIVS8Y8wF19phRRQB3eV5fAhxV8cIV97vF
cr1Evki4CTOGJQrYwhC4t1YfaSNgtGviNoC7IRVqZ1fz9R1T7x4cpZd6xNT8yJ6Q
WCLiNAP7jonaoodxWDU6UkQbcX+Zu9MXBwHADSgFq2CK2lz7mrXWoKWjp7AYLowC
+q7/VjjB/nwXg4yOHEXR1wo9Lj3/bTq5kbOPuxd8CmzVNaPS1jugGgX1W6CB1COr
9K6hDKyOHZXCKrqJWadHwE7mZLr4g1kDE2DiKyBgW13FkebjZqV+J2GFAACORH/5
wQiepyuDKqebAVQ6KcjKYo6Ytlo4Yxz0w+LNg7RkDx8fW3slx40yIreJrv+j9yCU
oCHPs4dgj+vyJyeVg4M/LchUa8P2MXsinZ2iQQMNnDPWOSUDJUBAH8xP1/eqL8GH
6kr7kXsl+Hrm4LmOw6ahD5egH++2Qo4hPXBbPACRxINeQEeGJUJ9LQa/hMWBo1Oa
ltb+Fv+nbl8afX3vPtwK3C2g9SXrS6hJ9/io0O48aepToY7Gg+A60vLiIgNzrc3D
uNOBkg8Qc3IBY7DWI/00q2ai46oQGTn05jEYL/Fdr04gIBH5V+E2UEHzdbck14Uy
IuJQlWpVdkrnaP0vrU2ObJdDL0gzpbLSZ3Z8v/DOv6pmqV4YaiNnsthAEWAq09gs
AF36dx7evRv5h//77ViXS8dC6EXuDqWyAEaWfL3zAfizUfHS/iWH3W8W9HI5otix
/KnPJCW88DuSL1VmR9gdxVVNENOQ9n4C0RthKWMpTh1mnf0hkdkTS7MGZq6PDAno
LrNiAZOjc+heaHpAulouyBIEpzqtkwgT70krDN0S6xcL64GZf8md91ZLDeKBSFGd
Vluk+ElK9C8SQ1FIzV1rTamh72jSQT3aE9K2UxqKT4GtM5oKaufz1RSQyCFXfs6+
V2iU5C5jS2jZHQvXZsKbk+KYL59h1dldA6t8fnULiIqC2zm4gEpHXxufXi68CvzR
FFzS5U+3YL6WiitPJyX84hC6Q9xJUN2rnLutiksQasWaUZHpZcD2WXnu+HJ5zajK
M1VSauT0f+8GbdQsDn1vtftgKPRx7J4NlM6CjwyWgYPqywwyKLQSkWxxnEkTq7yO
sI9dXwQshmA6WHke7z+Osmd1ai0REzGqOrCa0/uYucKEpG7ts2Iuh6ajXhPHGXz+
USk7AqQEDgMTBQdNxOj3Btw/Tw2CGLpblMJa1/Xwif3zsTJ1x7soz/tezrH651fo
w2fq2CvHc2HN9xpEPgGt5dHlepK0W3WirmsWq/KsW+jY95Tkv1Pnq7wU3OOS3KHg
+UamUB8AX7c/uQsG5CUZUh7MyOfOGToVSVGcYnHSqNJJiBRlxMs8YmlO2s3i9pC9
yOLOgIOSdLfNn+Uzu/Ny9d0xEQuRhHncbjYgxbF2pTMNTUHaYhp9reEv4jO4kl9M
KV4sM/exS7SrMF73ppJ/g9cGutpgXVwAf+xpZfQlXzf+/GMNduUH6JoY6RHoxW7k
3WSa831pchuikkP/Teciex+QyNsQv+JQX5sIHyZU6Uh8AWspCDiA2NgSRjkTM+zX
noSSfttGSM3BRV6QdxWAK0q7wTMMDokVoFGYnMRe6F6cwyDI//dKDqj0hAqBipQc
Mzc251Qr3Jevp7M3v54Bb/OaXfmwP4QEyY20RX0/qFNnnmUdO0REPVAUNhP612z1
yMSoAjWZwS7AX+VpqFDvFG7qaLNPjaJ7Mv7kb9wArbotNY3WoW9gPBJqMmfO1JyA
B+oCFdW3fekHVqB/oTS8Z7kURbzDEP2sNxtfG9v8SqSAJ/nuQh1oz75HqZNg0mj3
V+Q23uduOHgvyGkD75ciQN89b7NF4hjh03K8XeHr+vjODBJoG960T2b6QvXjNS24
RPtQW+GUzbE7e7asogBY9dBFq23wr/o54ZpsA2gRWDBwFfcjWPGQVIhwmyheK277
w26HIN1Obc77rykZvX58LjYaSHpN7/zwV9xWBadLMAGs+v8K6GUtLqIHbY9npZkC
vjx8I3Yi4U5i9EyIBr9k5VQx/+Zh7Wuj+Xwrv3T6DwJrGshyb4M0hOYIao1x4R3J
kzYK8T6rAHRvKRtEZmZMgh4zFFA5FLIj6EUn3OLl3mA1cJhWS3j783bIJyKcMS4+
5At0bWGWCdSMJjAYrq/ehFcWkpEA5OaFkxNC1lBLIxI28ub355u7X+XdR20r05J9
mp0bqWVhZ4K+4w51n1mAGLPrPunyz98eIz+ptBwQJgPv8Rf4xuAn4rHpNNzDFnA5
dQS9/wHHA5hhg1IVo7HMVmvBPAWJ1FF4fB8zLmVRReNRAiztxD8gJzDN69HTrH20
Fe7lw0QzUYWEXFyq1YjKooxSbgPldAc+5AA2Z7Ee8911BEwu1JkYK0tATe3pBKWX
1ePHzrn3/d4/afT99PGmYp/B/MBAUyugkMUN+qjcSQnejc2dIl2plxke1EOeuDpF
UwRNL2LhP0nXuiTNnVTMco570EK4e+skmhJjA/GCihuFuwza1nphzu0m6dZ/R5xT
oaTKE95yBPHFw/2p/9bn27DP6vagykTCXA7fyO/kpSaxtUuHKu58VTlevUk8J4GG
XAmKh6qLWvI9LnYFMA2R0eR5yLHRN8MM0eQBvJ4R4rDK12vmKWC3CD3XC7Yfq/wm
558A+foqSCtQ/lOKTsCti/tXXfKQaGiQBGnMnvV85u4AyczKllbgC4wgn6xvcAWE
ch5/JsVujgejNVDW5gI5KZYZoRGAH9TWes/t1zArqty16vlBEWp+4KJyP2zBO7bg
N4m/YfaIc0gBMUQ7ytSkOUMpolbFJz+iVOvrp3XO1T0rxVWMJPpcaW7kANQ1DYno
8M+hmjYvQ4SKbkrDfy8J4PIF+K3mUOfnItUzg/x2kQSqSbDgmozEeMGNT/gtQ8Ap
VlFBhkA5waEgHCPRS46/Dm8jjiqvf3z654DULVn+lDSpYtHQA+vkdAUtEhQGTy0f
llR4kb4afGtFPrWttWlF3byw4OdtAfRo06CBbeuUN3ChG5CgxsfBCHd6ILom2V/p
Jq9neE70irqw+6tW9Fm5/o0UgvSddSKmHj6C8QaULG1h5s8RAnO3aDx6RvUyve+4
YpUEv45uz2NlwR2OB2jRJxD0DYII//fKoqZFD2mX+qpVINU4dG9aLj/savEhSOQD
i7DuJUm0JCBAIVLTn8onXVpd73Os+8tKmKxhAYZO+SOeBwzSMdzsc7VeY9OUycfy
Qyzyo+G0gLKmSOqBBzimuwiUPHXJe/7bfHwOzBPo2OVYpl3mm82ioD+eIMQR8K2S
pd43vJrdIck5tpQ6nS9962lvv+6mJA4h9tV6joWwyZiiGD+SMxpsFviciwxUv+aV
alCal2P8M2t0nb5KGCVDKgoElommdCQ3O309iUwsibkuq6qOPD1zjoKJysELMBTz
Zq04GxlVsPQrPk1u0Uo+RDk0PJc+sIbZPuy9FLExyOzJsktKMDi8COnJFKDhz5oq
+dS4HBuCq9hyUW1ZjykEYzL6ERkHjCfITKaYbCix6+n0bxqYHPf6ey1j+AMgfMb/
jmgdhc7N+DT1kx+Dg7moNRzf4hDBPrf+5FpHjIDcNZwZij/Y6pdGNTcjbpb4Uacp
sycVt14LZ04KAD/7DC8TB4KWyjJnEgLYCwTPx383glygMW81sET5X6oMExhGeFPI
lRhVyfHJJdj74AzhRlzWMsw00ck3z7ohK6akhThzj6Krclz9nZhEaj0pD7XpOifY
u3DJq8ehm9FSiCAAzoMTzx32pEUdnSORfGGbqp7hM0YmgI018V3Ut29/OwVU73vD
CQO4Fxda0YZmUihwtAA9jVH1Z179CZ8L6rX5uT6Lb/UZpl3+qeDh8m+v6z9MSVhO
QcNsgpIEzznWy/QkAILg4Fx9Tr3z60YByK3/Sx+Eu7hXumogST405vA/F/noXBiA
aWw95U/mvC09kVfVre8so1imzEyzsGdrs+sAoGuioCqNJXGwwjHd8SKKpQZv/w9q
47n9eaA0ZqcCF56rk01+txxcocfb0T4ciSRXtF7RO1iFW4EAL7HaekLx7VAwmtoe
VdY+id87I660szE65obOU/I+ogJywgRbwvMb7fChrI631vbPmIgpYvWklPzL9Gxd
JUy7+jIbanpIzGAl+YD1ujdmC4R2B2WAzr35kVyC75N/2yt02h/gRjsZ5jEvN2yi
vrG/ACt0jlYjpcsNgP/4qC7pp9NqbHPONayQIqhHGUFkb7LIrkLS26IFPvrIUQX3
wbioQ50ilhSZbwmDrocEKYu1nyBZITEZ6839SLJhHevFmZyMtbz9JLyAPyK+990Y
h09eAY1TRpeVKWuU6rZVHIVMaJT+xiSfO+FWzFTGRg6Gt8No9ph2mJk96qD7e+0s
51amLhzjUAS8sMqHx40+c//WloUVeSqlVzVq9bf/HpCSFpRDshb3owTKWOWipg9t
K3blNRgReMK8ycNd8xLl4KBhusVdxDeNa9Urbndt0AtMDFSza7a9k1mkmqT4EvVO
werxl70skvtMskThXdikaCWTXecbX4UbAB4eV64D7v4GIFwe3PdXxKQL59Jxgw1Z
egturofQAkEamrDT9dwLR486ZhBXUNR6vxaYIXQXNAu3JJ69ZGt69zFJgr7C87Sc
FH+erMPJcU/mJ+xzubBsN+BtXDbNCo/qmSjtaECZnR1e7cehA1/nbLH/fax2MwTG
TF4VguWzZER+EayN2qaQwYtH41pZyfgNxxZeXNPDo7eqcf9ij97RemdfYcAmSu/6
LTg56aL2eGeDb51tdSo/vpL8yK5m95Hpyu0wHBrcRVr9G4t0K0HqAyGWNEByeHyJ
8X4/jY9wKABViZEKtk3ClggEmXBduoCnd0jAY6s4nfFNM/ybxVALjnDt9zWzXHaa
jZoygkyec8NnBPacbLLXY/xMVnwdCIEoH7Ro0S3rq6aQ6FiGmiDtdgAuyVpZlzmK
B/s6XmalfkcLjIKwxl0+vPCv0IFZ8mPkstx3O4+Sb+TmeokzryFIDXpM2vUaTN5S
edDUkp6Z4UcaXMCdAejSa/J5ZODDQl5+g3i1W7lWFyBOTgrrZ7MLrhZtHfp3cIlD
Odd0BSfiHA4ai5YNeBgUXYbGhd7MEn4t5/0J3xGc3rn2ny/WtczeEhPUfq3z5y/Q
MznuZ65wp1yICBU2Bd89MEhoHwWQuUm79VFQKJ2DpqbalnkqzVlGsAz4pL8Z7r1A
9Pomf/nK0Lz8EiBtZ44j+tfEdSKnUb96XeWg9OmAzqXBolo5OLTkJZAVpxbZf7/E
f7GgSKtIXR9dXHXd3VGlM0yo4jhCc8eMLUPate81/q06CBRKHxEJIGB1nJhdoWa9
N0n1HBvaATx3LrcLDtC/bKKmV8SGHxTC7rLmYagg5xSTKBX6uI945XtKt6m8keCH
Di8EZRVwq8ueIe5PJ55PDF+VAlxscElBSi6o5mmEBxr9RZ3iCd223wicJ3eQYtO3
5hJbrv9467IsL9NoFoo9/0xH8UnzDmjW+ylVUb5XDNeArI8EeCSKy04bKFvjYQ6c
aory+NoocX3KfcsSg4Qys7RJSkR9DW902w6GZMVqppZ1t9RUPtw2+/oJAOmURmra
t9X7DSqsYnWt3QQwjyvmaHqgbcfgXSGauXHDpwIABMJtSccqGsfRmtVS6E5VKnqg
zidiCoLC8qhQvsUse0OWKlbSxPB56ZGo1AFViuq9ACK7UJAwg21A9k8RqcxF/K5g
5GcmLPB0PDCIersVkEt83tZV+dKOI4suJp7r++0fV4qdw46tf8O3tHTdGAWqOGLC
5OFXy8oPqXLFE1byjTuOirsU07i6xKUOL71rzwjYbW7D0yvUKzp3rHeRxywaM+vf
ldeLZzkm786IBusLVItAqe3A8Vbnp2wVxSJz4ObEvozOzKnVvFjgb3wnK5f9ZhKB
vjRJvMnnIA86pTt7X11rF067pwPey7TTdOrFWIqOOd82jrqLdDBy9syw7b9jCfkL
W2zOkvQ4DtecZFgGZURFYs30ORUVkktP09/XWmbWT6GiZUKdwoygVj2BY4/0cXtv
htwFVuFOJT45trprMfY1NsfwyJwNfpKmj6caXn9JQ4BeVuPheAHaMGKv83ce0d9L
My5Zq0zeieQue16MgqpCDkHq18lFA9/eUs5B+ZE7AtiJcBRDik8d8+1BWtcRRCFP
nuVuAfI/Y8ZV0brl0jilONIRoIQVXX0cftdnC+zHh/XYOdlKzmKgn7yMlPT55vA7
4qWcCp2N7EQX8Q2CpES63myNuZc2vFjhnE5rhxDGdP1YrtLaJuYxjpTHhoAUoVdo
hEtEpznHoSz4WfrwiUXQYCGfXeoGiBo4Ef4W1SHSdvMPHb9n+0QtKB/CIr9UERZZ
3ivaXoZKuJUBouCFunWQjeTOH+dzZ/8vf1KEZBhxp/kqqOV6s8FrVr7f2klnMgV1
8CeaGLBsAe/12CQ3iaH3WWKqZjuiK0rsKEF+MyKUqz/2R+TaPO1rps9kfFujLLmX
zdiZL88gPuuGaVOOZABvbJC5zjHWrxnzatSHoq4i8E0cLvUGEygy6+wtBPsMVwIu
xDr5Cv+GbyhHqa9SZQRn/p7wGq1TpZM/TsoREoOW3YNhWB3RlmlGi4jToIAY/3Zu
ZUnMFG1ikheExIuXJM4wZF68N9UZjMaed+O/93Ek2SCSZ9JH0bAYxai+X8x+1LFn
4ZD+96+NNhARyCJGHdztRLSy+sFsJXATZvyswjjwWcEWjx3SXXnuCI9ZV4wDn6PQ
h+069agHFfg7QvmarznpMyrlk2xrlU5Vw5hp6hzkS465QWm+fkYpj2u9OyhGbOSB
26d1/bORnGOb1jIac7CJxFEeieNfAwq13grk/7wVJ3o6tbUja4uQwu33394J5Edt
9GtXm29SY8GfFiC9CCHCpfqzWTIcnkFZoWS8EvAUv4tcNMOAro2yENQvlq8YvuiG
lUZtnTHj+BEjhVaCb0JFTMO7APPXKh77a58GUo+eji33JtIpQGZ6Iy9lDMcOC84u
cNtYo0Jn1QwOqpl8bwdd5x4lvSTpndPEyaKk18zcFhTmF+j7YpwH2fyw94OSaNxe
7uwPFcY4xnY51uVe5e7NVbhDnvMov8P9+rEVreek+IWZNZ/+P5NblLugZi3SIYlG
DTEQ5vVfNmtE+2zFhUbBisc91dIDWwbOyxEvQDBUQV4mOrwQ/5u/5QG3mAbqIG6W
5Ql8bBoE2L0/vZwEFWV6VLHyTsfCC1RoUmFITNh0gZ9zXa+/pSj5UvXpuVVhsPOw
TUTiogftfpLo28wgHWqKMhURNGM8iGD3qCTUixZXWUxDGHwGdO7BAjHXXqoaKFrS
qmvv0Bww0h6gbOmKRVYPr4O755Hnobgu3XLdEtVnEt5eSZf3G9S80blcPfTdIuJV
VFUfT1WhsYoNqhyUniTaYwTKmcafjxLbD6MmoqISjujOHSr/wabf+KWU0evN/IWD
4iAOkKNsiOR4W/NrRGkXmHDxvIcX0twhehUwR3o5BmDO/gQbsvzQa/Z/TSofK2RK
yQ54sNNs6koDbpFrQ/8T76arstcZv5Knd9My8Ff6q0BeqCB0jXL5sCPn9pFWhVYl
WMHzIbbViaXt0BvEjVBAOPqW0eqLLbG1gmwvEWm+lroirhW5iZYDOKnupRV80LPD
o0CTk+W+Xe6vDv7pRZKEzDFGGMOlGEB5xE47jXkKF19G0KIv1QKHdEaYgBOZl3aR
xHuXGF/sJsIOK8hZLfN1tFn3KWl95y3MTP9u9b3mHQmrXY8lM+ylupkfbuOURxu2
jiyLT64rVrqJSEASfXx+AcZTRNgmAMqE7eLY/bvBn84jOgsre/0c0CUnWzpwtiLx
LJU+hwSaHJjjuPBBTj8krq0GDzJWxJz2YMFCtuzmY59kfyVmAubcGVevA/4vJlyH
tbYeJPLCEaMSBrPlbaamLgmmQeItPOkSUoK2V4OtL0cptSY/uniPx0CTYTV95zTQ
WRV3dd5jG0mUUMYT4DZqNiMcUfDRjdgZ7+qJV7EL3HnrKF9+R9QibQssONI9a1EK
T096BWZQH1zdyTe2AeYp6zmoBjbJNQZNmasG5+H8qUaY6EnK2EqV44kTJtUhq6d7
lUJAS1Uiw+e1p+TZ7VQMMIAjCFUN1XoaH3lXrbW7rKt62wSJvynHVNXZzmW7rhMw
f6kTFpCxw8iA+9qeMVUu+kbC+84bEeVHeGQNBzztSd/IvR/LiVWER+NN5PLXG0c4
SMhW01LJA0YbAYL4vXr6+38TZ1CwYSxP5YzxhyDWm8t6LfLO7KH1dLlcOS4Nm0Cy
aKmxoTaV2UlsT9Xmaf/NogMRE4pBQdP57ZkdF4jekDJ3H8ZT68zERySJyathmRJN
cCdHWAKRCqePL334YU8Cn3F09TQHKtkBgAMODyQAXBY6mxIcpBagveBXg8SK3Zmi
yWyV50iZYE3vYAL3L31N0/9m9gJQfislpR6WHzHSwI1BsboAp2iRklmarz2hcuXR
uf1szPKGZg3blDefopogpDHdiHrQoo8o7IK4sYGnNTuF3gAFtiNxyyJdlzyuoBMx
VRUhPIQuLOci0fFm2FODrZOa2HGPFvKl+N9dkOforAOyHdPrXoco47obqTQuxDEN
i4EMmRanJ2DsbAXm7o/RmOUsGkxgmofmAwHTJ7v6gcHTQD4RFaguoH1Wmg32wPTw
CHfsXeQ0hEVlp8gLJu1yKyFgYZkFHJKDdC4paMgAPmRCOliuH2DddMlAIiuuoey+
GOJT+EbGpjjHne8b4q0yVpREORLJMsOXMeqp+Dl0I3GOVuaW39CHcHjr2w2+Eo/O
6pcsTvJQzfbFxmjg15/H8b4EEweJlu0/+heq135I9hlkGUCuF/A/JqqfHD+hTEwq
ycLgVLBwr5c4+66l7Or5i8Qi8CynPKNjT7LFRVPn9k/XARD65FJvIxjMaOLD5xSv
HlOQKjA1haiLqXKPIRt5joKvVQ7Rybhmyfl7gSztP8+V4XJg8YF4//RijuZjN/pM
jdkZkFHxiqvBniD6qa+PUQbB//KX4/UboYig16KuIJxmGe9zFtjQMVR9QzqR9GP0
phBHMhJoGSU+6In4OvhKRTP4ALyUnATxRngPlcjTK7ETWjmlGt59lyozh8Go59DD
+JdgzMrc1IixAS7EucUVwsnGluh8mr2QmWhH7ZFFieKyurBSNK/NRphs1tiUtF/W
dVM7sswF2ScGJfsbheqRqICAxSwgu1wZrAkx7NpbCKgRzuI9nCT+H4TmDACM2uR8
ki4XkU3Ph3c/jQEDQJLf6o3JJopmd8N20BBK1cGZHlk9CwjKhPAjDUwkDZfZNYgA
NMC3Ru5bvg84JcpXMXWSym9MEfUWzwdASjOVvQicfns4746QqtgCkkQczGsiOlWy
A7/fF2O9dSRUaYzd9ZxV07+qYh/GrbBb1mEistXdnAtQLXtKoPpHE+Qbm/3sHg4a
9ibUP59rO2fDwUfwcV7DDrFVl6SXMSpz34IDdaDH95IXuZxJtQsoOnPfDllZvAZ2
yzKcTpsYyPOF9RFv3lguEZIPli9Wzd1Hkz/iLWIaY5Xs4KECXB7TGzOogFlWQssp
/JD8qag1n59FRkdbw1cI+4zY2Q7NsMmDn5AKC4QEuK0eF/dOWyygIjDTgldlkJ4w
lbLe66fMI9mQamH966j2f96IAsY66SziCzzPIxx/aBVqhGDo/ayfIIdP145OSv5j
VWuzuZqVdfMFiuFHZkhoVK496Om83QA0IB/dFJ7Jv0lkFO+80ECEUGfzXJ8ksD/J
028mp3drcU0a+jJ1IaxPjPl5pkR32yMUBNq51mMOQdFeWfoSaLRmZ8YeQYGz70zm
8IZNch6ElNa9IdQKZFrC8aivB/BMJFYh271K9uv2jy3UvEVScE85rtT7jZmfoYRa
ZYq1v8Mjc/j6NOj65yH0P6UQ71qWtbgFlHr/7kwCjMQvFD/1YI3Jy4KfCdAMFBC+
p9zHRUqqgHJ5qv6a09Q/U5drvnfp0lX1PmTW3JT9vWLasaiTvjwWxWYiAeLNQonM
6A1VLJB3qeWlXxtdqsiyY2ZCjVOu3et8H5M9DWusDz29PlH6anN2Wo6GV3jsQLTv
Q4rQLRh3o9+HRSdajlvRkFfiFoAE6th75K+PcfosSb6dD7VGyK2t0/EVHJMsie8J
MZDZCQ97ZA9/Tllzi9W+g4o5Nr7+LqCF8LUu6y5s1crhOz1Gz4UZVPVVjvpHqeRZ
ajQmSlS3H403+w6wBcvGlf+cBKXxsAh6cyXwCVZHxRdUtFU3TJhWuoKGQWw7daxJ
LUtJUuu8K+kxCWJqPepYgSeHTzsmT6XZS0RC/wdEZP2x/nnHOpe+DKr6vssGBqo1
+MncALAgbrqfcWPdVlb8U5dBTS8TLXFO38r44Grm+2Xgplc0PqdlxONFC62YT4FO
fmcA1GsRQa4JxIQmTV4FW0bGIG3qN2xW0p+IDrK771UgC9m5qsop7i4kkyGL33LS
DxE9l64Mv+AsA4n6IRdnmDTgpchi0wb2Oy712IEaJYw2UHwlPRDmtndes1/U+S6F
QG6UwHoz9gHvrKQ5gHF8KUz0K5qJsbWq8M6cXXfvJRGnNTrxOtGB2ZCM6VLUq2pR
374ZOD0eRR3phRnsIajAoQyBbr9lWKFyIi6YDKBBShHCRpPKk3VBPyrFFTgn+UBd
BNrhYpx95xJSwVsF9KjfwZ2cEcQi+AA7QzGZxasU82QaaH3DfUqguNKuFf+rg5hl
OLvdmENQ71pFVOrHPMgqLfUglZleOuT7UlxnA9Vy930iQjjTEnv/siGDN4dTXpgf
JkBZ7yePH+WhXNcOFaWBTF5dHtbn6A7V4aHvvi8guIB6D5Kg8ZGKddvtIqAp5tnX
MAzFAGqZ61/RrmDRuTI2wN43SLIn2VCfo2MRtYXe5OHqlsUMumxmIGjuXBPHAteR
5wJ0FHa0bwpijn1A1hEe2nr+nnLyL1uysude5Pd4Y3527HrljqlCLAu1sSGDNPbT
R8K58kaSM1cHwZGvJUa3nYVpUnM367lqn0ud7qw2h6bAqQVovE4nME6zG7JgRXW9
wORNsnsQ9UxAA9ugPIcLlaKJxmTs1bjfL6H4x9l5/abvN7dt1B9GuP6Lgd4q3xIr
UmFmbWrNeAnfv16ePnshRg+IvHFLKQM1H4zvRAemDkt5U9uU6QCYlRDmqB8An0pI
JbR+jn5LT3vzBDPaQCfmXPXmIp2vqLTUYEJNUKGDGjDp0r1oXDGbX1aslYBWpATj
OmzgFV8PXaHhEz1sdCO8dBQMAdQaUFfpxLzeQSv4be0ODHPhy5G7640/GVPn6sXR
QFTb730knlV79opm63YaKLhA+sLnEw5u3jEsgm/gLiG2wgEOq9nGYl3vgqntMvmZ
UQKsmNml/RjJUXOoOZ9ekeaK1dgoaWQSKWlW2ldiXH/M8hyF/kw1ax+eU0lMau6J
H/k20BnWbpn+DiJvHfuWrfDaHmdTtSxfzJpGgObuoVRpQh3c/ng7L6N93UynAs0/
3jS2X6mz59BQVi+zdXFaIdxyBejn3ZHVtzjG9O9+dum+3hJu3e+qiF0O8jWeZKOd
uZgE4gZf7gVURPndz0I0Zxt8K+iPWlnV8s15nOwiH9tfpwPvpJ8qElfkZZBIqgnH
ys9mu9qXDHgBoYHZhFEy5/beVXzyQ/OEsj2JfiXRBsN7aMZQORZJ5cciPN47CbZy
88j2s1kMXy+tKL84BkEaSPmS9ghntTHb+WME59pUGhT3mDCYYll0N6SNslONeEIs
H5pPc/hgjhJPm2XvdjyhkIHiB+tOggsmSkfnVowkVPm8+TIBfacZ7oDfBhV7UGr3
A86koQF3tTr3qSormz4RRegeTW8kbonxhcIRl8/xLqKX7bG887/v0P1F3fbpcB24
Ft/JqkIJec8uq6lscbvJgDzRaKISY4zHwv+BDvcc40edA+luYWBqRmk/CspSIX5j
qbOg2v1UdpRrNrL8FHi7UUhCggS/P4OQ2dWPI97ZjO7FnIaO2YBPc6sQcuwv4ltP
2Imb/sXiYJBm8mqu5qPRoYI+POWz2RxBPscEnZpMZysr5dWDQikW5ilJ7S6ejLu4
4Bp7yU5f00z2MZt4nXhNvY74pR8Z0108Y7dQ/DEHSP5WvpmZuFQfSwW0wffFAMUh
F8XkXqgUfSzZXXPYTW6Sx1Rm/UvE5Yv6YqUJuAxUgJXd2JlaAOzLFqfVsQjEGyee
ML1X1bBDF1afzIQ3MRY7sa0fJT6QRWUQ/6xFCwR0LPJrJzeDrU5GEvaWR2DNquf5
HrPXD1tg9hpZylfQIgVYVuaZhiiOMf/BJuea1p5EpEZNOXkGqb28rN+pfeZaDZN/
Kn7rjFsCZ4kWLWsulk4/eS+MmTtPwffXeCjbJUEuPFcm42mvufMhu0YHjti7cDXh
V7H3tcsXgGs8nK+PT80yakQP1N0JC1Ldn5qsNlWRZbOdI0ONLHV0DNonp87WecEX
751sjfRaFd05zWOBCDwemijsDylFfBeeoaFQTR/VSgWoR2OVUpJB7diQs6nhZuT9
WMt+7Dse1vvxhaZXVDnxCP8EAq2D8SbWfn3a1xwm4SCx2KJ/a9KNa0Jsb2Jv4L34
BPrJroHkTcR8LNqTEH4mFj60pgHAkTTzYkUs82wwV6iYNR3QhOK9whvJDfApxedX
cCT8k9ak2QJU0Hy1omAqLTJl5SGuygiy98EchDpW+1yxCH0quXdssdX+/t10rr5j
njFGyFUTKYk39dxTcRO+oKGGx2bjKXo+6Jirrz5Wp+JTKKlx+YdLesPlVyKtNITW
WhmqxtbdvhcuBH4kyjLWy/6l6WlXEv3BFPItFmkOrl7ow1XA7DKg/CyfuidLD9XK
q50XZpfDzMLqVHsYa2U3kvKrKh7c49uVc9s5JdjUXb1kfiuFBes++GEjO9DsoV8C
FQEoTyTvAxp4HVMRawRkQfv2AHJOjzDnqEGfBgi/i6mMjY86FHSJ7YAIgdSRZojY
KzVWHKtYhOdX4tOyz+8YI9JAYtWTXkGwyTjfkF79NrmKpGSqfTrOqLpDRx7bjsql
GtSC5gmx6BLaakFIcvibzXjjCV63RQyVR8//5XjrvFbkyxFjdfq4+IIkIAcjXiDf
C8TTMAJs47zeZXElk6zqpZnANeTx514zhfmVFEoVWeKuYG1VxcoIc298Xd1W0jn5
JAnO9iRwwyjbex0FmIGnQEM/ZS+Qe/b68JloUkMixVUNx0bvsc26VWGgnMLObz2t
vFOw6zJdVzNgIj+/L5jOHtzKlyueDFXiEj69F398ruWWujsv2daOZr3jAXFsDOUf
gd8HkkSLqutdJE9S0MgVYlXiKe5U/rF89DPSDav9uAUE0hAP9VjkFVDCZOXc3OcQ
mHI8Aaiywo7rhHZzQWjEFlLUXQjjp1gYVU70/u3qn9vgqE2i7LiOIH0yGj8V88XY
I72N/92gsVmvbn4kiHwDgQKYma+SfynBo4R6H7ulB89XaIwgfTp0D1LRWvL4l01S
CG2Ye1LQlM6gtCzED9S5mppBwTgWZOOMvkfUnoK8R/CQiDlOyaZ0g0eNqOWjK+KL
cXljxEKAXEcz5lb5kIQY7MG6DlttYewUml/rRdKHpmfoiBBfyqU1DPunLw2BGEle
5TEDFFBsj7UN53yx5PDLSwoNwr3/JKrr/Pwb2iADFDWqilf0C0kIsdUeAQMQaBbM
vaLLnIviqyePVhVzdC8FZsXunWmIorhMK8OVZkn7Vhu2iW4D/+MLg6nR6AtGXiGu
3YeigEU3xmjx/tPvGl9N1qTazlCTX9bduftq8IvYzBTu/yrCuHNM3BICQb5CDrKH
9hDw6c4YTvTBesPqRYYuHHkYMKlrDqHHBz+S7RzQDrRE8JaNDyqSVXVwRbnLX1Gu
ssuEnCA3ycnZ2SmbU8aUy2Bd8o6ddL//0ekJn1LQzWCwkWPkBybve5Q3v2R/1nmF
W6lwE5j+6xkeT9QJ/TGfZw6fBe4HzXk+ezgtovJAq5iwOtkaNzNMP7wz2jeY0MVK
MS/rGu0Sw/l8yeA9dYNeDWTZBan6+OpvVDILp6di8sJherSfQQLvMWLXTH141xrv
Z9aFt3XT/pZxDmCTWABYnudch+fbBBMJmb220mz5GLllWjDgEPkVE96bLPLe4vE3
2Webxd1O1ZzovztNIZukcj1cfMD3g+h0/t7nFWJnoRB5S3M4Ilo4BZF3syvf2v27
KdAFhwm+wbemv+uayeIZVBYzT+KPT0cQiQs2gLwpGI9mixpGyTvrAGBXSYpGnl6A
CGOl+F89flk6nXbu7Kmy+Hb/pjUjmKOFSvZZQsVRDSH99D/81H17ckFcpLz4kJha
IlqUkdcgjDWhKZn7LCdoSube0I4Et3kRvsznLPND8jurh/tMjqbiisjNP8s2D6tS
UhwsU5tbJocfJwv+fEjtjdo7xsslXdrmfeLolB0j71D9lIPI8V+lHfv8NHCRMPbj
+fBK9fZ4jNr8yr87D8BkfmfbI3SxoEb2OnmQsDWCN3fb0/6GZv9S+SqQe++0SNEf
mnbavfMC2eR/LVEhQGeQOhSGa26zy7LUOzetxtITLrp7kuFViLYV8VH2Ksyf2aN1
+55QlQADZHL3D780cpT/AjTmoYAR1XCeoZxac31MHZd0sBLcX5JvfeqQtLkhRPYe
WHt5DvdghloNEyN9SPC2U6VHKoyeBhz+2m8z1wiRif3od576ziCyVYSid8P+y+O0
aMjislGYLQM5F9z5LDtAhGux1fekZeASKI6ZJg9KISX5BH0q8Guelwmm9ebGmglX
OCmutYqKLzJafAt5uIed7KgaUM5orm0UiuK380feSetGjAd1LVvmeYUb0ZmqMYKI
0zQPV2r6DMxEuohX9KboIxXGYlQHdU25DTOv7kS0DTsARW4GNih4x3Fcpo9olX6e
75MbdLI2GcdU7dQY5X0FckcOOd4zRYuqz5bDMl9UlcAjMorArM+zv4tdJFhnGRCC
3YffMVBT8JTphF/fFlHeFUb+/ONgqxRlT/aaI6h8esQLkjW+E9dhrXmOzN1MQ3TR
WA41wPCfrjn/VdpWbDzsV4fg0MWKX8ulYROHL9G14AlygRS2YPu1omKoemeuqQty
xMEgjpiBg8JpdnvD3vK53NSEJjvLD11L/r7/86vZ5SEBMEfsRhSljiiaKtVVWm8Y
giWuOH1NgBHGOD+Oevrv/OCZTj2wfa3md1jqvHUDoYJp2+RTzizY8uEiPD53+6xJ
Fwl6g0mCO175lUQxHuS/5XkIlD3k7+b3pCuXXF8UFqc35m5spOWIag38e/JclVk+
jCrYBEbmIza5Ra0FSbVeSruzuqEV6vrmvFFByFeAK1vwLzo8fQ1ewIym3KvB54he
nCI9OxNmCn5paPjy2wl55JHA01jCp9+1Y/VUqJVhUGI1klklvWx5IoFhjYIi39Nm
dC9D/KucNFtKH3BjxrlksjnYBnFrj6JwEwVdFgwd6dzW4taqh9vSkvqu4mNRjLUI
+Hv5D2xbgOkjjmlyut/l3ERqVLmiqGvXyhmPPEka7s7wy2XV1B4TyNjkNQ2/n+kP
WivY0LtdheYRoKCv0Hsx6XatHRmlOTbnHv4g4X7knp+FkuwEwbSDmrRLDwJo968d
tUXElpYi+bAaGx5OmIc978TtERVHQ9mhLdlT32x30JjXH9Frno2FaCBwYqwCRV4A
USMC5DVn2PmWUa2lj7meT+CETT8RsPs5y90n8JOuuFvHe+quBPxSkAv//GxNIYDM
Fhh53PjZFus1IsVXWTkne/SHOIBWQR4FW96KsDLaqh6QETr8d7MOEg7FJrHMd0tj
B1Z3EhTO4wqRuhXkYWqIFhgn09L3yXQ+OeSeHr79kQNYQNIM7c5JZ5UgeVAzmbJ4
zmiXtvrbtrzbUklZ/ll7Q4Wza+eLtaEELe2+tuXtdy5DX9a3HkwUudU+Qdy3Nt6f
5dC9As4CMLalTSEnD8rm9fEi2DKJEQ0egZNlzVNgmr2Hq3aCbTS7M4xPjUsfc8Xa
H14ZCVNrt4agsSaxWP4pfL443IEGY806NWDYTrELvSw0h1a2DWKYOi51oqkJ7b2V
YE90iI1A+eyti2kiCdAsbi1UgxnMAupbaUN29nCuxjM4OHcMC7hZn7ql3AuXN0GU
a8U0AhRQUeO4LH7SyEBDo9Nt5ssV4CNxaWkdUvKCsOcpK7aJXHt5SQaikzDMa59l
15gpHhkcV8jXr/hzC2xhaIG7ylRkSrFEZcwTmdQYju+TkLA/MbKunMLqwo/Ap+ky
XNOy3xzBfjqAvFwRCME48scVwjhZJhUVDbIu7ENWk53jdmlv/CJA1wkHlomXMIrc
b6LoHc9g84i5c5ck21PN6esXPVKr9IOK/hZgrshVSs7Oh2zJqpcS0K3RHf5hRHVs
BmD53OJk9m2bMicHE/odUbZYMkrvlKEkv98htopwnv6gC/ECVW+dk9ndKmNkLW4J
zRd6fZMVjRs/9tSIXni51dSWaoUY/kr7k7derjhdyvsZ2f/DVUanFklF6EiYsp1e
xTPE3qBJICqs8HUbRGv2uSPGW4vTx7nuqyX1HTG1jP8BbW5ukIc41YH82xcDuTGt
2SgU9TrG3RUQPL6Zq9mgLcHAiDb8qek/4R/31neUL5aOVVdqMEvZyk8M+eHiBy1P
+HNqJvYHOz3RcA+HNNCT6yjTI0SdfWbWeCQfbO8dLs61ctLzh0OJjWM4aY5XhyFd
0EwicrcWUaw9p7GyXnHypdowlSNcXXTdaFLjjAWkY9ffFifRmr9SZzs9ht1kGKxZ
1LWVFbYqhUy/UkLuHd9w4TxMCztj3OLI1kJKWeZhBn0w9PmN2bsChUuTaKYNThAQ
LGCQZZMxcMe1TEyZeyny9g5wI1gerRe3gNHZlYh1Lzpm5b+n+YddFRV2gld85PH6
aXdcWhV69PTHEjvLqvd3I7O1oS3feoDSfIvM3tlv39W1l7t5q/2bkBDC+fKizH2C
Qb4nwgTfY+45oho3IWe4vMfdf0WLYvOX9P8/DaPLEOGJjcJRrlFnlVY2QpcpO2SL
Qw7+2aLdYsGp1E+IYV3eT93pV2Y7KTVTHRFTX/V2lq/EV6YZgWxDpcO14Pt+bWHr
hYDwDrA6FOa4jY+vN8lbOIWpQy446qlt4foEdublt29klqfikcK8YSbfLEAN9GtO
GDqC0DkdbP3ChNm1/jvrxcrglca7FQ+Ju3Ok7l89/3Mhsebkln3ovW7d/fsE++6s
FPH8QQijDJ0Sbml9G+hdw+fd+2orLi3eXnDl3i9q2csZgO10FQcoTGHkr54UwWxK
t6Mj5ohiqM83+KuNKOt66o0a0uFbtTw2/vTU+aBE/zfRtF6cJzzJnTTNWH8mXm7E
8QHJ4t/OpH0KeMg+ajx4O/YQ0uNekyRMOKEUFtl/5LBrSZVqsbf7hVr/fyAuar0q
iDTiX8noyRbnE1yO7jYGw8B/e5flMrHfKtPK3RFxrnIzOOGkTVbtnnQkV840LC67
IKTMm/euqUxVFEPRaPGX1T8Ugk/8YwF2l9rs93eszHNpNVvZ3xjPcjecA15x39ll
CBwlRyVo4VTvP5e4OElO1YeHJz9YDXPVNlOhjAj+ya2xeqkabKsBMUPp74GnrhYz
oEnLMPtXsB5/V9JWF84Y4GGd1mFLEYbd6QjKemqZqSE7Agtsq4qvVX8gq2iUpMZj
rzFJRZxvq4bHMVdIk/2RDsu565YDD00XO6C+dhddahOf6hParfPFisR0rMSFeefb
BliR5l1i1E0Laxr5SC70KNbRaIdI5ZDiUeWLsmzyuKGsM6d/YODo4cS+NkLYncwa
QAfcKR2wJRzzpEVzI1YUFelN++3PW5NublFlgK9PRng2RU3r6oq/k5MsUl6XOCz+
GeXr64jg9Aq1cvWrTFMg+u3zjMdQpi5HZibubPrmjJwJgjNzDcfDkyGNPM0HWl+c
JoJjMEryZQwZpecONbt5kLXFnwBgw01F74CaVIubCC6JFShuAOQJxyZ68bfINvN3
YL3SgB2SBOm/OPiRDDzTtMtTdXssOZs8KiSp8na1XaH9oXQelmw2NXglMywgY7Ko
eHZQKqD8PUn4TjpcUJje/ObUaortQm4ZsPyVQX6O+Sxpto7AWdikvePPHkhWuo99
MqRdvgv7HYrJB7UKKc//+tw05/BXIoKR3iu1ZSTr31GyZHNjKJIuYvrwpVy5NRyG
ZDPIYAo5EMfEya8odbrezrLzN4uup10BVP8P2cmkLrbID1PWmNoETKlC6WXerkgs
G4wO0r87yKOZXd8kpUiZ/yq8fgQJPfZnPYgNWI+EOb9ObGPFSYaxFwIP6UIfCy8i
zNjRWdAVV25OL57aT8Wk7WIN8Ks3Ft49jHv1RsDBRob+GjBlEOund/MZ4srveusA
b+tIkPvcFejUaQtV5DgnVeYSH17890Uy//o3fncsL6Uh3A+jmc+NKBvq0jXrd7va
EIJGwBx1YfZgDJlOHG1OOlcm2u7qeeYzvzidnvhg0iBBR/YgPPvzBUdzRwTP5TI4
ydNudlYkAdtEHGZMa9o0OTtGWRvD6AI+N2LySPT5PRc0DqFwgBgSJ0rArNSy7CXn
NgCq4nIotA5nsyqw37vjpodBr30RzmQRLww6o0zduN2XDiK7cIiXSRIuhzBgNmus
TSn7V93PQb0O2nX1vNo/nRdCTzomYO3c522aAcAxxU8HRQ1sKGqmySHq1pf93FjV
A5ujmOUE6aULG5e9xB3esKPxaC/QZrrfffkhWZ65eJi/yX7oJTF7B/wx8gOonTZH
4B+aQuPsx95LEESkx15SArt4I5yRiAKvE1HehE5KNZAlbGIeich7DMUxZXQFLU1/
8vpbmXNLVRv7BKZIOxdKO4eJxxym5eOuxpdZuSUBq+O0RuV276e2znq+XZ03BqIj
L7r3UZXHhRseEi3AUFD/c6cwwkKeZDGl8VQIHlwreKsnevtsqw+qiN6BnKe4dHwU
VeJ9RvGug7kt0oQihQxpLGN8xQBzQdz4Rh7uM6jDABTnG1HVO59wIY+sUT1/GCKH
GVHXg9PadKGlTPZ0XX98FcPtFcdaPiZ9XuM3zoOantWXlENmnPshXVz2mbgq6vPU
lnUTzq0Fcz4eFjrhFo4kIPJsP7EVct6po9OtuNLZclF28Hx/s9h5XCB3U7Ds/bpO
GVIOupBGSnyNgwQmyiaDHe0MRKMKxJMVFefYaFGPwMJcy5ZbK/oRqjvHiJtcN6Oo
COp7DKfevWu2FZ/wCZIR+kLzjEToqtRV7vAZgDpqvpa0deHhjpT8GAdYGt1yiB0a
kQRvukDu7uxYv3vnWYkMu/sqcqbZNSzvE0w4bFn+T61xgWzDeXecpZ3hvsWd7ju1
VnKWcB2MXbqYKmnzDYkgqwY+OC9cmTy9qAbLvZSW6TMgoQP0FzpGDhnHzFEmwDKr
ZY87QKbCExoWGeajZ2KsPtz7t6wOPn/E8mL2/x1Z/ZOiDKcF1j1LIvLYYC6F/AVs
le99yjEGNTJfRoEtzP+CIG+KrVZ80Bouy4EvMZWic8yAPdJ5tmblIEwPo/iyjd6v
wpeaR9N2itJAt3Y9Z5CDuwCjTn0eMkmLOh1ylxHHxa247pVj1cNGWp3Opq6aXUYE
0t09e03pw2vUghOkQODaS6onoTAGB4SuXR06NwbNXhzd41TzmnlWiLz58hPWBS7d
NtYprQqXb0mcrbqTUOYh4ZIzXaOkEVoIjqsVIwcELyGg6G7e5kFe7ohQltckeWSq
5PFygbeyVE9+yvS6NEIEzQlJXT/Ln2RCoK9vvw+iGOouLzUjejQVpNqi8NlOdtHX
igFlDUzDuCEkXNFBzanvX/L6hYZfZWAPv4qr6/LKfWMuA+EPxUIaOqUIb4F8p6OQ
9Rd1Lk+FgA7RHNoMsnxPS2roxCYNEwTjMVDvTI47S1xL6uxDwPFRHLobZeSQ3QjI
Li40lLNbPosDhUNadHYUDmjYxENoAXJeN4q1Tqgh3kdP0+qEd+cmXkiNF2W0nbdi
2hRCqJ7RD7q52vutOIqEPFWgbu0vkYng5DwmV9PdcwkEcv715ykdRgerHOHu1bbr
axArJ/gljaVCA+2yDrWa+/lKKzXYHKq/OH8HTKLrqyckLioluI2ia9sUeGAomZXg
bMJlXOpCr8PbhTFsMbUNM+0Rl2KW03Jzhrrofq2cJFlgQGA4/Dn/aciQF+HXVvpr
EVMQf+9zne3J3/J3A1Vee7K8r2OdHWmGWX2OpUyY3Ck3iIZEXz185irIZqS6J3KY
K3UgYgyOgOEaoiOJ1ZViis7nGUBbO/cQE3ikhRvFs5T33rjmIm6IRGecoDL1Rt5t
YHYFlSN68XPiGUyyz6UyWchNz6CAhu/3hwEAmZJwWDUCR5uMEI23QTrAUq25SBLm
QE6WITlg9LGPJVaa8QS9xtIkB/3zU05dLts81XcxtMOqyf3hiuuZ2Q6CwfKW9HxY
4eMrVf6dUc8XNj39YWVa8WZXgt0bZdjE81NJaHZham3JbljEJ5pBKb9+E0087EkI
QKV+Z65UBmL4UfrYhrDfHM6T+SOS13nX0EKKBhGDOzx8+Mu80ZKIyfMZZX55m57A
+BeJS71az1THAPcbw/hg3o3+4pewTH6qc1VSXPSjVOrW4rn+M64PPalVYOkzmZ2b
2GLS51GUjsb1hV0aZ+WxjOQiu0WNUNdkU4v0eTEH0AN2Jp/8lr3VTGVKQLdrIxwW
PnotqlhNCTLWRt2AkDOJF/kplxa/+VrDXUta4/8XMOxFbXb5mY1pNRTQS6KpfhIg
T25gA71tiVeImmYJDI/9abPyjlGyvPMG3kisTs8GSSdiY9Ahi2AuDO0ssdyRkUQ6
HboSTbioO1LRsToodSooV1Sj/UmI/IRIbYiRurzn7ctr+LbMuGFMbRQo9HIXF7UP
yHbEn4A91u3ApJuZ9pHTFNGEdhE5ambg9fKMGVv2l3bfiU3cU2uM1CDnXlOvlh4Z
LvKSsKiFOnw2izCaQ4f1Rh8YUYlzkv1IpcJNMAp0pMPQpRcv5T3WCOeUS69bzqa9
4crJmiCtHVFi5EDt/rfBgLJe00T2iBO8XzgWM0mtSvEyeV2gKiPhlpNKkfIp7iym
1lotvnVrjstJat4i7ntAcHenBywvvUE5khCYvdGQNJy82pXOUk/foRrCb7T4o1+h
DqBfzNK21tRrPlhRmOPBQG3iOijIlo51x5l/zwznFMUX2N0HV0xCAV6/drBRNyVO
JqpepWxOy1NVBD5LlK8XtIjbzkmCbNJEVgHLJt58Q2s2LcTzLoedvxFAK/i83iUE
NdDY40wZN4g1lWSfridRUr5qwh2KkYrzf0RJwAaZxsAf14O2jurmAeMuZXTxC2Up
1b9KxmPpG6OdVwsSlT3CQ9KhiovQ1rRNz3mMWB4YW6vDigZ5Assb+CGSGNMr17Hg
UQtOOCnQviHfzyRsjzzpdUOMTowCExCfZmvm7U52sCUwXqDuU2vuZp9PGCz1tPoU
Xww4Mvb8huX/uCGbSrkSvWAxwuKFvq2ECbDvHpDaFsSwbeqZFMeqFUyTPg4tDC4e
P8Qzo5bzZrzaZ9/2Fam7oaRDavrktbijtV0+dXbum20HyJe060f1DodwZR4H/9HE
0tX5DTmoR/R4e0SdnpU+cXPQkdUEHqaupwVh8yR9/t1KZ0RjW2L5837jRDitQI82
Qku1aH7jEmMyWkoeIZ0HTjnyIcnJOUBU7aiZONpdWBDwdcytCPLX1H4vnUw9Tqbt
bfSz5xm/EQhBRkprbykfSgBxzDO9lSkNDzzo45w5vz2fEjAdF+PQUgrjbqBuFfRQ
O0FYJxZdsWtCSrlNkd8EjjZtMDSjB4TR2sjlAj8U3UlvhtYtFNGHWVcf7VsbtTc8
PXLvrq1A3tlbRzODPmaeuZCwD5cCj5hJArOKQIVUD5WZaedtD9+galAZUFWXVWp/
MKnt86H71XOyV/9F0CZDGqs2ehl0jyakiYC0h4X4SG2El0knFNZ1Dy4f/zbD5KXk
ZFbOusU8CadsHQlEfEY72btKDe8xCSf08qxZWELqwZFd8tqmgVmm2+3A4ymRJuJi
IdNuNCmpDfbE1lo+KclqTx9Do2+73hk34IZZIpto1OpFcmfVd+b+JdAHHpKgF8re
mszNKmkSzyDTXr78k/PoDrxPF7a0EXIbzX9P+8D3jGqHSMaVX8jMHtNHoYrwzeAz
kCSqYjp+yAIT/JYZvI4/qE02MmpDCw1AHxxNMOAQ5lb19SsQTZdvXoTW+YLaKLdP
U7MdtNsOSExoH3tVxXY8jEqx9nBP8PW68sVm1KJWET6wlbxRPxucZRpatqcYAeIi
Rw41cmAgopkAHie3QQvVOWkhmKVvXls8aXykRHRePXCD1xZI6Qh5W/q5nIarq5qA
nFTuxPhpsmfvbeCIfGUlM+dyINJ2pLVhn4OWJwdklMsyaY7QEWs8dTtkjznwZM+1
XVEtw4msR3+Lj+XtUah5H1HgMg1hkF1QIJw4g1YWJiFt01TjHQDTcUn837WRwXOq
mK4fhUaPNncp7H1ve85K542rCAf/nD2Tm21QLsvg8XteHNLbzYQc7KI24w4biHJ6
X0bWO4i6C8aBuKoWdcfe8ZH53fPLb/L22gal5ef8KIXs5v2tsFOP/DIWDQjGFjF/
0yITJ8lUwlhkKBBOtjBmUQOAffigYW5C4ekbM76AdgV+IRNhTbCgfW4caJw0TkQ5
NZw5nePklz7Kef0Glh/ifzW8T1w60vRuzUyVGCLJGsCAAZPrYIDNWNvdtS1rxy0Y
tPovIeGMU5ltq7o48EsvtAIhq2hW9cgTjuABd5NfHu/EQDShtCFWPw6+yTgAu32m
9ESGaWI3/TFgcej7f/5HIGrC9cFiYVWM6V8e6kn0VTB7lGpyAwer0+Oa9kvGVAKF
SMTUustSJC5biTUtXI0z0WEALD7RB4OH6Kzq21Q4DpIFYpmLAJ4H4YMl5NTGZahR
HwNl9LxfZPM4IcimKXvQt1CgHETeKNtzpsvcqa+qThLD++pvVPL/KjZ5VGBQOHTQ
UTssWrZ2FuAqqbcIDjTUnTFv4BN7pXnNyY69/pl+jxZz1IS85eUqDi7cDWUUch2B
vrL5VWk7D9pwlQzTlx5MASm7tbYvwt/Ahdlv2cluQgNIkmmWlnRPywmhznrbDG0W
TuyF6zr8hHH3Z4uZGQTBEd96EtqID+QrfBu3gwxIz0ndY/J0KAtva/ooIqjzHJi+
PlfNQXWmFugpIysplxhGd9t31nCi7x8q6aehZ69WnY2ZZ+m63AYw7QL7PbZa+E9t
XXwE4VCvIqMeleGBcvM0bPDlMRAdTaRXztZHPqAirGL1VXYabhi/SQD9XUrFEybe
vY9X/gJsTXv70Gh8MfhyUA7pzxJxWB7o6IeMQCruKpgsy6VdYVCPwSW/BKwWgyl8
i2AFJKx/trlgKUHkpK2m+JqrRrERp05cJDjPhtoG3Hz94m4o/q8uSYyB/n1uRwUj
tg4gvW01I2GSWJju2E2C3DdHaE2FV/ddDwY+TGENnyfxkhxmMTTqATU76BQ587pZ
EQW5Y6h0UN6Mqee6aZ2W3R9bHlR0pSyIhrpIYWS6klnOlM20P0gdRYevkj7r7IAO
2OOPFfIFGMeoKOkrp0NY5r4MSkQLO0iTyWeZSn/j1HRjzTQMc03QJKhd4JcIeFsx
28CIJUBpVFZYPAq5KqoWI5JveGgZGsWu2cfcg+YJJLTuabCPEdSWeIZsn2RMabcc
NTD6ZggV/yRPLRKO+DmCe/r/5ufB84ZVxHvXOEkTcD5bEVVwjjGT8nSLF/WSdjdK
GbQ0E3Mc0JZ2AfbABASk6nuRIPjacnFnaNOf93EZAg2UNScL3QL4UtYZQyKarvH3
bN20f3+TNGw+2P6P/NzvvTDze+WD8tquk5QbM7oieZaR8zuAhtyhOEShHsFzi8Qm
g4f/hGDLTfTTKHuEQRh6kzrGVQhT8gy18SyWDEFukvOrsbKjwcuH4dTSaOOzZXpp
qfaWDZw6/efx3V9LdMv/IsUu2Ff1tXL0jPntEOx9v9nKlQmU5/F9Obv8bELpFfgs
D4PmGJ5i6bsh6wgHz42Nbv8oiHglkDWlvQbWGxIgM4nfDqj4E6l3ASS+Dk7cgySX
w/Tnb3wTfS0DR0PZl4J4o7Vo6E5mdt7jyZ+PtsPEBZVLxMigO8S89t3ttna2JjUD
TaiQt5EWVUxBw4L4nkjkSgcOdnVCqbY6stN5hhVis/wybniEB8WNehyeWg03AYI3
2bQbzzUvjT+I1w24UBL5vmFAmopXMv1DBBlARvwqT+jIA8bMRqbhQ6PoIeLxgQGu
q8nCyVG/EK5PDtRT2K70wGCvxRtf/VMzvPuGCnPG6fjvA4wNfcZva4xgeMflgabV
x3E21Su2BZ3jXLadZ23fFyB7i8siOlcbz2pYOZJyT2QYDeakKIHpxtS7eRCCDtQM
qlAR5rOjaVuUZMkwMY5gLqrHVEGKeCQ1a9g4y17Ij+438NF1KOCnd6L+3R6CLKcA
r5VkT6c+f55mCklIXx/DB8p8y3NzuEU3icUsUpwtSgaQMSHhnRW7KZHV+tSYj726
Qz5y18OGO3TAEOri75XEfvCiKh3ncJpT5f5Qkgyk4xpMZMXYzqQfZR11FI/9UqcK
uRm7917dOLfBnh3zY2BtL491b8Z/PJv+vwMHeLKKH9YwJWsuB75Ca2ttetAqIz6v
gZT76JSbVYS2V8x9dAEOzQp9iKbLD2B76hKblqaJgH4YqPwuGTwiG2bVgB+BfK2I
6F7nnW4u652PSx2QyC+hsgyWYe6pDExcFGfKHDgURod5XN/yuDqpC1uAxY0kCdJt
jvwcR265b8PGqdNQG+g5bzoZJGfhDLuVMb4myxhlSozSXWzlVUVhhZmALUWVfVs9
iMU4uZ1weObwIeitAwI0EqVT/t9R8FZ66dhP1dYPrc5rYsCq8+X3wBDHEVhrcAPm
KqnTXG7+PhFG9GTbNE55QbcuLO6jTBdnxMVntlSJK+aJP0dlNyX4bLN0wmQo/g5A
OYQjJKdIAmw496Mwcv5wETAq091zIReRCYNMzxGNU3MAFef2eHt+No74Jb667FgJ
7wpffsSBbd7oAiQHLcqRku0eTu/xoOCdKCY64lmk0dAlgzqrxM9PR2BRV0laUvQO
ZM+/9lk9mxRb3ydMIpvP0LbcuNI4GbTPSrijY1UWyxkexHqoxXBV6IqvVqt2XOkN
aBijoAy3rEMXxV9aODQOZbZz43mwe77+7QQ3FpJv0QDz761jfZ8s93ACkv9x28CR
CGLXY91Qlcqm4Ep7+QFzyxI4bxfm167pg4/gI9uzzV8X/J586+1Eol2RgJUE4l4E
OgxrSvDMAGAeLRtB6uwreyH4Lo8xFHZLY8UBQosEjiUR7B7/yNDYgEIUGlC9xa0s
X4FuP/DfUJGB5UdBhHiR3EPNvs8vzFszOJaONesdc+oprIOdjLfUZdyeiHUJ+4Td
3CrxWCNv5XuaI1pOhXKwtJ/ZpQIEUSOWv+k5mOp5BaFh0GtfnQeOh55JDsznB6z5
iRCgT9wTHTpv5ML1AP7PoPZQ6L7N5sDzF98QY1xLSGs8s5NDFzGlKaIQfQmQn8mj
RAFi3x9Ppi6WVEUKyPLLvwbJU/ScLB5mrWhDlUjIiANuIStmcut0kyib8lwiSTq/
v0itQluM8Rgesn4VRDglPRlseORhKDdXupaRrqCTp9HHLHmIbYoXmUmbiLB4jMAk
rFGWv2qWeA/+63RboiJf13Wav0LwWR9F/WbfzGJkjTXX0/KVbYYnGdhTuqCvhhS1
ZMcnst/GOjfZilJeCI3VL3e6q0wjLVmWW70FsDgsYtyb/SCGT9IVDSy9aLO2nOmQ
7Fswka/qJqqANfbd9G6H6jVc3PRP4ciuLuIGfP+LodJI7Px1W08DTTGFF9+zSGna
bQEXQYulNvBF86bfKbv85oL9sqtAF4kTgI+dM8gMRHHCOPxHLdWXRWQdzoGia3Jl
m9sg9tVOQulFEDzHJ295UrjOVupKD55INmIKK0gExoTBkSQwfbxjRlLBr4xhMavM
4svI1DjOY5H8wbCW+nIMnREBC0b7t5ToONRPVZXHvLk7XJ5E8uNtKVWkQyL4IMgH
yYVSpjmi2qRdEQ+vez/SP0KZQzaGNQ51ZuvWjkgoBRf7kKZY+D2ooC3HKhLsJCdA
qEa4erK4me8KgnB3AcI3FdOvYXiqV52XChD72p/kk0O8KCAa1KcJZWjxHO60BFO6
b/Uuyaj4bKrWSRFUPRV9fG+rbvHVNhLPmepluCnu+TWGVnLWrz16MNvxp3fRlGEl
Izy2WOioIvmCQas+dj031jHLvwEO9mHoroqonpVbte5+esGqwXlCXE6KCeznBHXu
H/Vw8x1hyIA87/AwGhXXCM5tsxfEMnXFq/qsys9md4zWapOSEv0EDdV1xLDcR0wR
0lnSc+dVr0QSDF8b9aY9DTyAOxgcdhRUgvZCmetW7pFmNjyXF40+h4SSdhzGft04
GaFstzxHgOlTJlK2wNwcPD/Lp/B/F663H42B1HSHRyJLFdYejpVi+PZ9fboC8Ukm
NUN0p0zIWLmTCaKHMwe+ie/ftP0IENcgeMg49JSaemEpa4s6OzaQ/3ot7Uk46/CK
hHAZ3nh9O2DzdYe0igRm8HEqfkBi+PntmXocDXSm8fLRkXdq133FSrxhCY4vurl7
t9YM8p3+Z/FnJOopmGKBK+7K5NMkFxrTY3LgBvsz4nOUCm6ubx9FVo6iqqGHbknW
xgYbwyieyPpr3we3hVEft8z4cvcjeUZw88+YtHhgPe5ejwsp/EvudKaKld6GV4zE
QHt7WSeAs3J0M78xuAAr7Ido56gR27g1TIZvEgLCH9oJfNBJpA9CYJzVB7R9OYlp
woGw7O1XnZ5xn4BxhL1KlSjOJ6P7dfQPF0w69j5AD5WwUNbVrnx7k7ZDw9dYTiL0
J3W2xGkUftFF1TbR/YCoO1YYv0zhvMoxOQ6+l12AFWBprlZsHMyUDLyqCMGEt/E9
uqQVxNwMD9tVA/jpaA5RReBY6Va60U8hzpIHBK4jmi3PwVANN8CN3lMctXn2XJrw
A4JHCpllHc/jTEbRmaTdMEQO+oZFQkTUU36wgjVkbCI2PAfboETJpcqsUjSssYYQ
dZStl0F6+l0DFDWydTGg6c1iToKYpPcD5fVmo1hEK6+WVOKzd9bx4zzLZyeRMoWl
HwIB1rCw+J5wI5k0znkQjR+Pj7+Fx6uSeNFkDk8TX03x5gh4urH93QVQBP7eoDPV
BKyrxBinjQHNF3KOD0Onzo5AOobXWKuj8SkApWXrlK7d1VG6nYC77TxeW3lrF4mE
blQZlbJTVZgVrU4Pgme9LaazqzVL+42ZXpGPp3nHpSBlXCqTwhXimn+IkN5doBdb
aXeLwx3ncHK8xxBuelubLUlEbXvM6TcMsFezcPfoVHD+6WcfkxOFbje69MBB9FFr
VNAjJvHlHJB7fnFcZrLaHhe1SjjVmOJ9MTB0jH7DA9DE6WgYfaURppi63fh0SRQc
4utGJawkTSHboPmkvqk2m7toK9ova4E6pL3QhTUxmLobiVUs7fdFUZFN3nRM7j+f
VxJUG1JOx+TqjdfT1ZvNMzPpAUoKysJBpRC8cY2m7SOxbNaTWR21aTNufSIsdZLL
L/WB4eAc7mEkV8s4jHRwMZijfllw3V8vrlm03vYdqd97SPcpzPJQnYJW2UUwmUfi
aIlRfZqa9YGG9g2d1MqgwhcQUjunhC2naGkjQ2YB94S/iNKYKS5qI0u4OJrhPdFd
K8vKSDJnohLDMvujcVW9D0Ha8ksW9XZBx6NxRfKgGC5SULEqHbBSE8CsDKA5+LqW
y7+qQQVvw9HLWAE/ua5uFn3vo59zyCO9d0xraZvb856+WVeq+5MsDF0yCN87aWG5
6oQUlITzc1Tnxza3UwnRHttCa24Xacx6lUH8vVjOzCAj43biDxclj7W/LHhCqAst
0ya886jFjakFC7CSEZx0Qr8Ragl1SR66EE53VQnLVJyeo+hL96kfmj8shEgQSclb
enN65o8HvLU9fjWIoNeqvRYXi5Gki56dxtedOc2aPyED4KBt4ZXkSXVhiAyZUEyE
OMNaOdYoROBuATWDC6e+j0PHYGjC1V+bhTHlA4a8UblD5/REZ6oWlVXNLqQFRXzi
6rbTTLMemVHThqcoyO/QWYgDdawZ+OFD6+XuYCjr6aYdYDJZgfbQSEyxh0C/PgNp
RqPs4UjEDL6sDPYRk+VtE4SmrhKnNyssQL+j7K4qoy8Gebjq3QS54oxU0jMmA+0J
FISfawCDd384z2UVvWysl6UwlQ2ugw7peWY2WlhSIYWN7r93BbYPaogBqlgfCPRX
dRbBjcDeplCtvh0RW+MuPuqb15LFQay0lA7qyPljXqGZr538yFWeUDVjKrXzgmCb
CXL6VqkIpQPmvrXB0C6wNO5EfsrtgXcr6i3/fjXmBZ3TxMWvrOvY2KB1xIbWv492
WZVOWbkHIvOam9FNefBA4UhDoOq9A/uNRCPOn+coizITX8TwM4nFnN0+kkAdf0lm
N4yqFddu1HLVBqs4Kz8hxXvbvan4tByAinrsFEt/pYu8oHv+0eRShPjvmL4blbWI
L1ACNvnJhFtwqj+1TLvztj30TdRWI5Z1thiHbk2CEvCpn6BVVisZfWKshfqQdCJt
Um5IdvL27ZEhVWp+EMtKW5H6NRQjz4Zj1/NzqC6fhUlNT+rIDtA5Nm3tFMUiEVmS
ZD/3g0lsL/41Hri4uIOj7/YKwmOebRuHdS/DJeVYmOhzMS66/cACxU+Uuv4Jqbim
BKtjZy/kRc0rmrA9rvGTrK7/9+jd4y3roJL3ocOsxPAtRb2gLTOZVzzeRmbIX7Di
Sqkzmlt22FrPXYdd/Qin+6RGuONKTfAOFJrh0Oh9CQJPW5o+ckvwZRZYe+LU8ftq
7DRFM+f2DGw/f4bXXRuLmlO3qXovDgpWPmY0MM2n2ZZM/yM0Zi2GwWaiRaKP7z+x
4gpUh3NW1B2WeHZoHSV9Lm5HxTkBlOe6H1JvLjuKp0+mClzr5pN6+rQk0wYjfqB1
sLPWIV7dtapd2nVpzfJCLEpg54MmBTdlufJMcE6LVNQJJ0PbXFh11ROiCi82Qu7W
ZfKVNLM7mxyeItckCgPpyMKbJtS8IXFXO0bvY6gTliljE/of2hczu/dnWoExKvn4
Atr+ePivOPcXxlrUUR8JiTE0dUK12+3VZUWNxkSY+7fCxNByh6KIT3m58Sw9YvNU
CQEaLd9M3GkL/WuXP1RtGOxHssmykzI/vS3NgyE6r57Dwh66stA660b1iwNhfBDr
UlLWFR0a3iRgczdHOtWDGOQDXmC2VUQewb/VcEw3HjhpNYfxA7nVizIi4KMQXO7B
KJEJJGpIxYEZ3exxiLBWAuT13sAqyEmL44THdoqtXoJ0CZypynJ5AbdRW7+/XFfj
Ce6bVWvDaqqA4l5IIQ5zreRKLSiTtUIC7mHwEoj/Nc3oFKY2lOuBMoe0UtTxWPfF
ZX1VWL5Oi0fbeMShGKHqCff76udOyA17ROC/A2DfAFqxpDIlvwLkg7w66onqXUrN
khzwBULVM3zXjv28k5/gIYBGZO9Ly092gl4H24yqyRIRJv81eF+4SP/Jn99DOILw
NpJsEsRrisqmJ60Osv8mYKs2TNr/TUNh56Tf/vNzLZkFZ7A4lFbzNpx7IxEjAlsp
z0s6hs++PlBuj7yhfAr/3uNht14j3hVOAeG4GJ748V/vQJTXL92uNuaD4oe8KH2X
lePTZ5YW2Icy1rxWXzl1JiIng5M9hcDeHqdFmibf0KLwPGtmwkhG5bbqtSaJsD0R
ltPGwZ2H34YNQrqmnSImx4ZDd0IMiMs0eLFnfsPjsRl71IDtYkdrqg770IaOVG8B
xyUePZK9yydOx3fXVSz0ErWZm8Uj+1I4++pwnAs7EqSDjoMnF041IAASiogBSljj
IySNAWpRkUjwPjaGlgy2GnIFG49w4fMAH+4gZgziOmmn5z1usYdmSoXkOeMUIWQI
aNpEGXrRf1tOySfyfdMf/LLlIbJnv2GX4dWfjnbhoGcpqxBtfPr5UpyUxwGYrmem
zFFpqfnjRf/DhsIMsp3val4MYCs7GF9rSo6Pwtk10Rk6vtCwfLQTYZrsAqp+LrBU
DXn2Fu2nlhoABwpqnDRgcj3l47uRLxwZLL5L3PW4mNIIajgMzCaTbiWcgb6zXWkX
ilqDsBGQmdiO7ctac/4fkt9fO4Fia0pTYteCwlQukpInkFr8Y48XW08OnN6CMGPU
Fg5btQuhi2dF/oln8MpY7YxpcrW1RwF3rX+Cdp5iMlCGM4v/FHHor0ngFY2soRXS
CG1jLG+pOeR5W//px+j7oh6FUzjUBlulul0Beo1o5Iu+TVaDXpiqz5Qi6iR84vDQ
CsOTEtNQ8N4lwXK9mg/Q8pDiIk6rmNcKBdMgTXXOUNhkDaB7GTa6NfST3+C9aoOb
6ciAdejQ2qw6SVEk4Juk5NnSRYNbYgQvQLf21KUc/eKLeiRX5a4TFxcc0hIW1l7Y
6qFgUYbhapkFrUGPXUJ7JtYpTFUEns2KNGyQkaUDHAYO8noGP4zQLoa0inPYE4eS
IaCKfvRzfxk/DvmsMelCxpq6rHzwVCT6Qtq6WbYta7ECVb9BzWOejvpdtowTa6M+
zJOmicE7kMgul/QcD5pcwvM17RrkKicSeznrT6pvwRncOHd0r4vEh+E0G6hlSKNU
TpdUuSpShHUT/hJ7/XauE3rFGr68LId1oqZhvwC208KX/XyhMg09WyzkVOPWvjAX
PL3sFvdZGlZ/ppb54K9Gum0ZwxnhIla5XTkdccDoS8W6mVb+xbaQDwIhBD/ZMHDF
bwrMSJS0DU+7fors+zonEHv2xQVVH7id29VvF4//yt6N660YP8En89PfUdB7Bpp8
nySj/oUIMxJfhKExCGJA4bax0SfBwpqStFR2DmLKZ/AgcOjHSm6tcfbbAPwm6uYd
efOHJet007aThuj/c2nxCiUaCLx3druxGCXCTsVlrFralgYCCEIVssd4yHQWLp+Y
MjvTm8oBnKyjK5dQxKm5+ODddgJp67NAbKx+y4dG0E4iXlReaTXT3vzCRWQYPqg1
bXw27VXfBoJsJpj9UKKY7L2es4W2Z8nihMvjxL+RO6fZiHGcmFql0SFM2XE+sG5E
1fEV62HDE4y61ac8Vycfg0lY3K9d85aAjX9Dp4xUffXZOLoNdJN52tUGh0FZafu8
5pJ9ueV8tog62MdXisOS/VkLpdVS23JDcOAMfHJStkz0EjaYEhCV2iewFgEtG42q
9DBLyubFRZEJ3MOlEOphdCTKllovp0Iq6B5qd5eeSg9L3GPq21paFhDHKFJk+C3K
bgDyozi9R0ilEABFLMEa8wFTVX2OalAZcaA4wFUQeamR4UZyvF9F07ALH1uuR2Op
7u6HSLaWQld/dhsdIX83O3KaDNyKmT8p597oFQzuCNjXeUtwRZSyflWIIPJr7FZ8
e9otEh/vvKcr1o9Q5ui7oCA0/ZyuFzHpcePay7OTryEzbFjG4OnoLoZxzUkjPqhz
IIPqH3v73UQB5ig5u6J5B3CmNvplINgswmvQaFGuy5xk5hS3RkjmF83jvnYrP0dZ
EC28zNkYL6uPQ28QJ60iZfBTTBb2+uB+QXD1/8QuVlpUMhD6bvwFnXQSbB+mfGrH
Re1Go+XZveYpuNRDz1YS58unnO9adwv/D30GLsCzJ63rYPe6Cd1TUPNetomb5qFV
3mxbI2NCOtZpkt6rjhctP6fOGSM+oWV41LU7jnEQXQhAXVlLETC62ymTm/eTP1ro
u7cer+0pBwjNjIUMua29h/BkSK2SL5Brz+tkcx9ZQB1Yg3BLZ+vnzrOyN8xBcAVw
KBe5HoJnQd1LAxSSn+9O3+MpIqrPIVaBFJ50R3zS2M/ceL4uyA+s4ZmTBvN6Zqil
iC0sDTcTeS4Px/jeO6Ejxrsx/viBEhQtPOC4wHW/ULdyDP6RfvinfAbdLRNE7Dkj
V0MDaa+UpZyZkXA2Rra3tNREjo3EglaVo7zygVJB29LpcrsD99GtTINWEmjzUmmI
XWjQNsw4CeXK8qJLg05kT6ngSPr7pVkpNEoqw2I1x51CdBusbb0pF8HUIchTM1ru
Qse5L8vOp4WOo3VcDSnI7FNcyYlclJZyQ769XUVeS/UHJ6zwpKrSEEWiaK1E6TC4
yVo3JJJV3K/D/62A7pbCLZ0q87rW/JYy8oLYxDN5tF7p81D8+I3xN2QRRyCVYmeW
t70oqS8PYvyfkPIMicBZgmqmaRyyq7gAX1X7GVe3lX6qY5deEi1JR8mJbynEXIMA
maizH8kSwfgm0lzDk+UfAuNTENk6R8DPMaOO4VEiJbD1su8H4iiF+yubnfRFuRhf
X6Ap8+RIWFKg9vP6HMs6TMLFlJwgFMItpgNEDpU42C6zprU/4yB7yreJYdDZ4Kdr
7weuZiXMwhkZK92L/VIcHb+q0fIbdZnx+Djv/gZMmE2grrYDe3aH5/zk08VQpyO5
vBS+QQ/AvDbM4mNppvb91WAJX6LcAb1efrnSxDTFnz7U7bDIbmiCV4igtGbQUdIL
DR1akhRYBHd3N9x6RmQoGXtoxSoGqwM6KbVyoJr4UybYq5DUG54JM1nr9aFatV7d
lLsj1sKFAAf9nnrnelPRrTaRm4bvgPEEjUx7UB0Ty17InDx/XqisLBSCPWMUhiJg
soREFTQeKPuYnu0lmu7XF5dq3zC7P2UrBh/+ElccHjOqGdL8cSxEkQFTfVqiPZ3/
hAozE95CL8cTDFzE6yw7u0DjAqoQry62b4G/BLY/j/5chtptFPKRF3g5+lTG765+
dIgKFZkQFvzojBlXH9fj5wjRNw2RRI57Ir0BwRC9DqiX+kpwmiQLW8Aa0W/ZL8BW
mzF6XW3IN+rRhcG01OYtbc25wjxAtv9zXQz4q1FJEHiKZs1IDGvul5CSbXArnSAF
prhpDxWL8cWM+UNd8bvMK+7iz5Bw2VXhyVZKhBhF6xQSzMTIZEEpXqn6zk3DeV++
Jjr/VYNeebwrPvVlsUgeFTPxesFDDJjDo8jOs4aTUfpyYi1cyiVK3PE9SRl0sbzH
5zyKQASeau3EJFK3Cha54Dg44/UTKG/Q3ueelt5tteWbH3C5mK4evxiPZe3k/sXc
zq+i3y9/mLRpMENuoG/NlsZdsGDvy4aGSQpwivCn5/gQHc+SiNlwHd5dnM1SfXu7
K93fEpwWWxjKOM5M/xCN8naNLhoN/mZ+0Nkbw9wnIobL2XmMEYdHaXroVsrwiWYb
wNTWY6B1/t1idthMWiBI7zzlyjKOca7C5oVmdrOSVP3WwaXeA/cFRXgvmucLkWkl
H0QEJi4zrSCjdtM4/JZfEWEjSlwrI/by7BVYzcpOMFQGzZujpfmlWzQ/BeG8yCVZ
2w+Mll57Oc8NlQR4Jhd50YonxWTZJGgphHarAtVBIfr+M9u0PWaQHEPVjl2KE26F
YIsv1CRWfAJZdJgnhsnYY+LZqrYOG0v/QvaeA9r/h0PwLwMhATNQMuoUhJSkrgmz
RXswsPBnCMe0+Q2qSjNkqtBgnudk+M+qe/eld8vNmhYiSBoy9wmI9WFxSuqHxZ5v
+GGPruCBHGArFE+n81jK5wpr2k67PZABXdzDKEBfCYg+I6E2H/MB1Ywp/hDGgGba
aRvrbfUL88Oc67h0nxO/ByD2vTYEx7RUTbiN4Z5oDfwv6WOnD3Cl6lsu/jFGaVdz
lBG6RCS45k0b9W1gYW0c9fC4XIkFebZaBfQso4aFSf5bupJVYeQ/VcLrjkFuBNHL
WCSdUs6h9XZCWDUWtWOJ6mKzF4eWFnwLD4oV8JCPG3FcUa6lXXSCYmoJvQJv+Mzi
V8fR92xrKxjBGcZpKYqmzDvYusxnR92FbHXPnAD0KkZqhrWQI+SbJ0Q8jEQXymXE
Kelay8rbU8Zl+OKtzEmIR5/R/zBwsmvoBhtOCIqEQbX6eztTSxXka+4Bj9/Fw4wg
3+EcmhqDvJP55U4No9Kov7dsVd6bQClvnr3KcR70LUM/vupVJbIFHfb9D81WRq0o
u+rOaQ117QH7L7V0ksKl36do1SUwnigDByC6og8AcYfM4xo0t2TZwT1woaDNCPnp
wVyDxKaJtJoLqTflhgjyFW2VM5vDim6cjmbBKaSR35Gw0YGHsdS1Ayi3K/bv1uH+
z771ouZv0Q8tVAyKe+FZs/mlEA+PANm+Vhp95EAoPfNzUSnF69VW/I0FefkibOts
c/WKwxEZksDfkhpmLBWbbyjyuI9Z86O8KMkadz79yFqrCMsspppys+tKQ65hesM4
Yx7Z43oHurP/EQq0IPUFuEz5QWGv66XuTt0vtH2wp5hrvoBwpikjf9IGIs8rRC/A
BEWHrL+zRbrDyh0JmjENUIH2PjlSk3EbiiSGlsPViIjByXQMgtdvgiQoEXq9PgdK
xyjhMy0UCEfyD45FMJw5KEPzqJ9cZm2xPAjIO4o1xRW3vNwiKUzFEetPlo+K32aX
BkXLKhRjiD8v3BXQwsFad8pI7YHuDf5B+vksSAuwY3Khehg1POl6sM6vgtWQqzPH
ePfdgl2H1kXQAaVcKUqEAZPdX64zZQC0cI9a/3x2cGEyhf+TcftQMbEYuwpGyeqB
k3IcbFGANc2N9QIb1sDmwcz1bHgCXPUnPQOYbuSiJ1sxl1vgt2/a4Swd2KVIVoqx
rhnUovwqTWsG/psHFzw/TK11KZbHE+lJCyzhzQo3UyaXpc1jvbkUs7oQzytGZfGv
poAhcXVJM2TawC3Hf32QNXt1BICJFYdE5xuUeRNawjpcMPZstpXnfm34zY1Yn9Ce
qJWGTmTLszwn38H13rrZ3mNMjkR7aSfQKahuGg8PR5+0UapptChjSaMi4yv9johl
X6ldHcMJ5Jh/BSEy7raKu/z/XG77KctVrPk4zIils9mt2W0LkZdIAZ6vKw4eVqIt
bW1x+yd3bfLGSMWT5J4mgWW6Gb1VFYnoRoL2gPciCfB6Cih83+aRhM+1B7iC5G0Q
/TS91Ghob229eytPi2IJI3QH4ujmZRfppPQa4oWB8R7wVfxLzoUj5HJCFL9JbtrK
6idofggLYLpFj2HJpgx1KNfUwGJ+otzcHyEjsvSbso/heW43zy44+mTFp7H2Y4cn
SuwvX1RhURJXlGC5/t1lKQ+eiCnMfxPb/ltB/VoFFbPsqsZmaQSW8WDnrnIGUhmr
bSKyruu4JrUVGlFHVsSWpQg/O1THr2gzJKDFHmNdV0deZxx6benr1VggGbTiWZHA
aFF7vuWpieXMar/U08S6kpBHgktmXmLQXFyU2CquQvmNLAQ79Ab7f+AX71gedmn3
OAzgNKF7XnENCd9m8OP5P33+4VdJ84TmRGZUWO+4L7DzojKFvSRY5q1GYv4zMsnP
uqk5tgXJ3cnFjvmTIlNhVCcsjPsp/IFUdyhh6sq+E1Tm9nldprarj7lsPWvx51U5
nz5k2A8vYE99+ZH3yKkjfZhcVVsbX5cbMq8z0km8zYU9vfJGXdop1S7YsB2x3Ds7
/z1P7D2qvHpm+bUXQemKSbM8cgff0zP3UpHBorVAtwHq2sdjOCwR2Y7bziB4vlE3
T6iOe3vT6XnuCH4iynKcHP81Kl6HuVHc/Yf/Nfvlbhq/iFYe5xrGSd9IooRiqnhD
brFAcXyhltlnT2U33nm2adUslMnqUcDWeGU/ipRAigd0lh/1skNx3QFKJOPzy4y4
zXeYMWwZrin29hfSpmx7AuWOrAnDNmu/VzQxXKEQj6J+m4lOmo/cuay2fYJ1MhmY
81sauiNteIGgyr6oedRCepzqE5tCW+yAPdsJv//bMeScuoCWUR9AvcI4ELtU/mwS
+Rgz218DBugJNQ+HeT9KYbaJ/4Ehb5AfPlMKqrE/mMFqeR6cusb5I2Melyw/O1Gp
nmw3/L/jjmQl8/pUB43ZstVkCWficnE5vcDwiyHStSZ2ULreTHx5kw+DBarc+738
L7GeJPvXwAD+gYmmnsp2G+Sa7l8dUVS1Wd/FzcRbwFx0g6WdBxt+QUE65Fw2MTIh
+yjb5JzQIxnwL/CaM2g+j03D3R29AKAk49cmLbtDzr9t2EpbSi5xCREVMDyRxJcm
IV6N6rO1pWoMobZARU/yXcl2MHlIrIhupNVD4SFiL1MYLVtyAtWyzwUcLleNoD7j
lI6w7PTjK/EXavlpzYCQBmD8SeL1I4j/guJUTgKateQtj3bSlFO1VpDRA7jmSnjC
tnKX786kDhxwV5VxxGoGpZgYLSRO5KmDsIssN2hqMPpSHX7RaWGOxekixYPG7eFR
c0bg3hovj0FpR/aKN1FUlvrru8ag0EEx5KxnnXcMF2/ulL60O9P2iUpzS/lMRh4y
NdEoGgwVZc/aAHcLCpUwq0qMK7pbQZN4GcfCP+SNR63EpbJPtQQV8W5C+/yolnzz
CM44tOJ0sXAVOqxHq42i75TDYGTGHAYx1vcK8sszY55y2CBPuVFzNucuwwXOEorq
gRwnQUxZ6qNs/3GCs6bfRdD7BqizAHKm7eNJQPy1fzGiNfwcFi/C3Eh0zaefWRd4
0Fs5ntzqLTRk+Bsyp9W5yc7djqj4u+fBnv31m2h9tXvhDS7o6f8hr1TzmaPOLaVZ
M7zaO7hf+zkJnHnaHYr2FVdhkCHhwY29vSqID15qqngou6chF2Jo0Bb38U36KHl4
CENr83Xc/elksaXxWWEDhZVpkvsET0gNQWB+lXDOt0L5OPJuqHhS1uVTO/3II7M0
gbKIegJ0BaNPWJ/g3Ye/e1IDwtQvhuraBp9WPBYFC+88mqqoOc1CB0hrxEKZRe/N
0I/lrX+DbqRpgtvD+hliqqPgJOjOXPJr1arHTjRaAQRUaN/FIpLKjlJEXHPQs2Ok
HETRecQz3QPTxnbWNldQ22ql9k2nxmBBKGU213sYm/p97UJan6MFwnZa0vOJJ/YR
XF3py+LcfTZE/Ba6RJ4Mur5+Vfk6aa3JJ76qAXBvhteuqBquFCQPMSkXgJcNCQX4
VeTEUR5t3PZWfoOm+6JyJ3ABvCyJi1I+b7d0zQW1F35Jj70mobUXt7djbOj9XxWn
WIfEy1EGlu3fT/D8iFos7lVMt14gxUHVd01ZMlQtwVDwx2LlyvHKkyiHgGLMtkRA
V5S5OunVeLW+RnECE1dmDYTYL5aS76XswzcFnq/Dc+78cRMVngEGZVQYM15TzYo+
ipG6cV20xg+0I4ZNK9W29qyahW6h5w0ngWm2DLaRjiwh7nayeLSKYlssD2jY5/j/
PQmJvhW14RRD8DGYmaYVFTDwq6+t1GxLbBbWiFpnERoZUGyK26mKxcxPFxvlVxLr
Vlr3AJeWBNXpGq87Vh7YTovAobEnnTd6PbG5V3n2pMe8+XLfuDI8vPilhhWdTup8
eGPvrBAGinw8+CLkOngEYcjsFfuB1dRrQWLp5SsZO0XJlt4Peig5eq33efuC4WBl
rJGoaj75bZPX+cjPD0TShUrBle1+YbKHk9GfpSsT42R5Ldl4Zc3fxCyzbVpnhhtz
ac88LlKVHAZJYAIgTAbuJCN1wZ1vT4qDYOQk84kUVtfc7/ZcyzfJItjyHL+M8NiN
Xh/1+5Q3n9g6qwDcV9XNIc+uDhDOoFjfJ2k9JacTATxaYjuwX7u9uTYOA0YbzUXm
RNdf/mbSu5CyguFKjETl9yT5V9jzuB8aPSISDMXVxc9D/SL7VQssheCkoRqYYv3d
Cd3SqzzL9qI4Ol6Chm3J4k6c5SxmqVbG9zwGbMJh0EW0O6kyQ2DDIGaNRvl/YF6/
bV/GRbZlwdf6h93ftZH/1tr3lcgaE5GHDS+Q5/cgTDliyg8qsJOkvyfZCwYmeCQg
f36OmUcB3FaXfTkW7750Rxs7svGqjNnKf8ttBapR3EUzxi+h1UAJ+PyozovwBpol
B5VdqxMszspT6aA33OaRahe1vBx6ZRJoJERh/K1WQleTFVWlwkdpwC0XMMHGl0ss
g7COy7lZvUHvgnJcYZml2kfYStcM0MCRYuk1oRoqJFGHorXPe7qjMMmbXtbKFiqw
KckD1ZLXVxWjNo0y8hfr539mAL/ioUQhnIMf2IbOgB0oY3kmbWhKYtTVa3EGD6bv
liMu0AEt7eJbvdomWBf7i7KOW8uNZfA6TtHKJ372ZhfD/ViS+4/+ny3bykT6idUy
s18Nq9UBDA5BgGp3otLTb5crU3Q5MNQ4F+1zdmf7fcBqMXQ8+7tbdD7uQ1l797i2
Ssbwz0AwP8eMpgbZG9IEfGqsJ+erB9rOIFJpJ1V6mV4Lwwuz268PUGl0UmYB+3to
Zxisnts9BDHFbFwGhjnYcG2tFv9IoDZzVH2T/aCKQstLq0KWSDvM+lH82Yq9VZie
pDfECbr0rEzSERpgSjtOo+nKQaKENww0R261TzuIPEtCnxtN777heITpDw4MquJm
apS4Cwkxm2+xMkrnIZvEK+Bx4dMoZ2KLWMs6G0V3jx5ZEXIjOIjcGg1ahyU3cvyE
ye23TVQ7nvpp0pEx/gat5A/K65/jvl9XIP72F0FaLt0zLccwO6ta8w3KKAYHzdJF
rQlEvtwUZXKPcSnKgeV/2i/rHA/81j9uLkx8SPD5W7WcDWxbV2Gh/GOkhMtbc8DS
qu7nVIUN/F5adTKwmEVL9qdqPCjbM34asltFOzZDOqn+AO7CzZhpWrhcmGE0oF3e
7Oc2b6+zviHC6muZxYm/kibxCoAf1Y8mOl5t+RTaTNABR4cedvRp4hkkxwytH7GW
o31MIZF5ueyTgocqSlwtn43vSYqyEkQ2t4N1GG3myUZNq8OBgneudTWK4/4b91e6
y2pWV9vCasTXRyX+7EUm+/nYvZ59OCwPo9GAZcHOz9gBhtU1wLGaYa7LgCPWsQD0
S1vvxrTD3jP8rwLhgx99lB5aHeUMN2z9x2PiRRrH2JMEswmtdumvK/rGHT8CB0TA
kkmPd0egLsDVWShtOyss/zNFSuievsyUupq8BA39pqGldwevwuM9IST5uPnALHX5
P22JUbvBlSjCtOLUG/MfwRwwVngs0kdXyG181jtbqPS3Q9QgCNyhdgAotrSdIx7P
3Ve/0QK5X+5hRCMhk8r3e47nZj0pmmXAPcEE/w8krEXxVJi0ZexpwCJhIf5Pi83x
c6RH36HE2e3KtScAugw+84FFT4d6OrsJul6JHmZ1y0FN5QyflU+4rSNrU8yx0MlA
1jUBJlZTcYfeKfkUs4+PyHmm8SUvNFfgv1P9aarFD6TbApcFWNCRmP3IvnA0gBn2
V4m2XeEFfUEGzgrU5BVeYJ/XtEP0lpQpRCHzM90cPEIE1DMono5/SfoMPW1SkqLU
vW2PA8Ldr79kFk8jLDU0q8bOwCdoojjeVSwDPWwSkJcxALy1/QPddAOdjP3w6IfG
Dde1EcYL6cdr7EJIwxMkq/KEDvoXBOV9+y0kjrn/fGmYq/frzvABKXvN4NB0SXCP
hpfCW0kdXfWgbpWBxaIaFg9NbikxyAjFcUckdB88Haum+nYugQ4ktfZq+mZSIOTb
1x3WQMxRp53x+jvs6AiXL4UMaJG4vhcjsBKARZeERi1tEjChMblZ7oeE6jNzlmJx
+Xnhp50AZqToRtxsryGpummpX+5pygmSgwPy4jH1BVe4PI+D/YuPAcyTA8ppIt3B
sPszslJPQIVXoDj3iGPAN0H+IsYwtAEuy8h3BrR5smmiQVItOPJxHB1llrbKqOz8
p/xk8ZwMeeio7ZdFyNSuPYQLXjEgIJ52NKGDY6P1hu6rIkej3qSSv6l2ftQwCxTK
44/uLUJ7T4Nu+abP+V+2dE1xj2J6obt5d23UV7e/9ky0PGYypyu5DBL7LCupsD2/
wWoNTszqEON+Du6/5IHQ1rESVGr0HoPLOS7+er8r4z8QI7JpWbi5Cg9HHLfb3la8
d1hEWEam9jQW+bpT9vvMu+shuQq27TCJJo70aQs/aN2qvaYhZytPtukiPcbtV/lL
su2aITR92LOIoKYKH6lOBudB+qnpnLdGPK6Xlv/TE5RjNmH7ngMgaWldJhgJw36J
u8sk6W69UVRePPppIosltrQa3Hr1tROgNMzg9M/5wLDwMpGqS1EIi/s/mFvqAMdP
62bLb4lAx2w2wx0HBhIvTcFP8OvDfd+bohj6lw/SmE235KLJE8DxpWxm3TGimO3A
p36dvH/BadgJpk+cRxTOrLYbrjwPpD35HIDR6PkewXujXcARjbPU3R0tmjDI7VT/
ModLtf/8Ceeunhq11opEZbOwinpUWRBMxrTlClyHElwqbdDf3fCFineFQVo4Ll5T
Ok+ONbTW5c+ZdPw6YIQ539tkDl0vw401qK8imL7t3D/DLI7ahThN24ApkDdGCCs2
dbzY991OAheDhPCl/sE+Su2NsB7cmOyimaSBREKtTO5DZui7RmO0hotuOl+sqE4B
lHhl3n/ytuQhKQGY5SHxXTLtw3QhlU7t+gBfvoEr5exrkQllC1J+ZzfxvLz7yfmt
iqKHZ2D0ooZpVM0tuS0oa35yJSof5DNsXtSt+dp4r6B3Yg66B/X+XElaD43ZPT0E
JWvzUKFb3hRWHqQJXWdW7+lG9yyLh4APxKB2M0ba5IOa1j/bXy4NFY77JtwOFJAv
cRz39ArHPkrX7Bvm4OVlN6VzBKsye7W0gZI1Es85hpzIsk0ZtsiJ1vBnQkKYrOw1
PGMNbdYaUTEzhhQtLtm1DrAU2ayamUp75wugW5jQN1pLOO586XDo2cwNtmdSWCBO
YK9rYoz0fwAZ7iRWVJBCUYCcKI5xWfLKlTaY/J8xNR1wWiD6MpPxhehXFhHQkLpM
13XR7ACYu6Ai2F/um/DDRjgREGVgN/Phu165O35ccY1l3EE3DFKIr+O3tV7JyEtq
kCF77snGGkXrdTTAgJ0En/G9la0pUFrp1YxukMEZ/ZRjz78+FmQXuMbn6/n/qbsB
epj9s+cbya5EeeoHT1419e9MqIi7FylAwZZH8pCtDooQF9mgOw/xpuhH/g2/ROua
KQ1CWnhsJoE06e5imojWbH4m4hpwUmDl0WnOS0D80rtlIgdw/HH1OIyRCVZmbqId
aJWC6rcU7KYKTTi1IhHlNAYoJCmag8dCiigK0fuOnV9sKlI/UJ82eL5tPUB/RYHK
GIrau5ui7gx4wxn1Qq0pOeGqZCoU9DFARwZ32yYEJMNtkubdMxT9UE6EyycLzGMU
KP9sk5n9dKENovWCpZPPmnAezTAP1feV48rG1uBnPMGBjpNr5tEaI9q+tCGpRH0N
3vvoKGmO936YN8gLo4JFBqjKkhqgdZ3MKmnKSn63NNr80um1YMKj8iJAmxgur8mg
N+Jpo/nv8t9T2RomWbq/dIyRNUAfYGyKNWHlQkvP0GaWeTQwAioeaUEjtimyYDsn
1m71FMirmTzsdmUfFcjL75w6kpT98xD/9s0c91xBXtnTPyTQObV0luvhG5W7Qh8Z
Qjn8U8vLFvjNsQ+ujid8T6GcLPS9lJJ0yN9O19Nong0bA+GQ0K/Tqw7eVox3JYTj
Tgrd8FvQ8670zcoHFEOxRZLalewQvGba1pBgI7sKzduNzwy80RNgIUYcmxSRuAlg
pisRPKVaQkWAitWI/o6deeC18Twl23DE49KMLg3HSZbYs2ZHJm6BIKRxDyK5T+iQ
vVncfGn6HInd+95hGd4dKa2OKr3oy+U1ZSvLTp3k5l095zxNeap6D0SjIvvVRGrD
BK+M/v7AfoPHGLSQhbKTEwWYkxrjpPMy8fIFkYbDYLY1nR6oZPHPm8uv5TeoMPmu
ASpfEORQu8ngb3uzwbV9Tuct5X8egWWCVHcJT2NstSHRXsl+aK5nVaAEZVTcd1vF
shUKwi2wOeWIawAgcgP0OotxH2AL/9NzbqZH+To3aqw6IjOBsHzjZjxnyd+HsYks
JPeZKbtsGedfPMq0ZetsGQc1ho3KDL4jkD2043ApxMuHhgE6wN5XUNPFx8Dl+Ncf
kDaHzd1hQpD+UTnwn9w3X3APPWLkgK6krlcQjmKTtuLPByRm4C6QZAh41ZmHJblG
CjFPZ0NEaMhB4PnA6JOAotKOAqIokpxHW6KPg3S7wlNi5GtMM0/fUAphhbPhBbdl
xToqBk65Qo5di2TRhzEDJIciVWX5GmFZ3TYPKLxa8J/20cECt7UkH7o/JymXZMx/
BsLNOsVJboOrfU5BImzVBCIf8yGTFCR7e1gVpeJFbHtedz1S37NbueGUr8vuYNWc
UeLmjHFabHjE6pxKnN7JMIWHOpHiNwCvPlx1kxvN9QKMv1u6cVuaclls6GpCIVNL
Q9Ne9SzeHjMmlq0rDluQeihj4O2lLqYERXacfHxyu9V7C0PTM7rOwDim0jw9b9bZ
JRwN5CRWlBUZJIehVwmy2XHZ/1yMgPDhRtqkKr/cev6vRRnHTbExQsgYL5AngNvD
f7irYIChx1rAQ/a1/2Uk1cl82mOlui5q7I+NsA7DLFFmsvxWXKfhYL585CnWfxok
dEQeKSsPCFjEeWxR7fr6SW3mc8kUiWXNibM43vD3jreS/vp7bMhoYyxR9b8Jt2LT
UI0lUHWUarfxiV/qW4u5sbc/tDA9UQxfJ2gicX1ObpGJKNqrav0T8w7om8J+lO5I
F6nbkuG46hTLAUOQMZwMPuFKY7qo+Jyd1OO9eXTK72T7mizfGz0iJLOf0FIG8Ruu
ouevw81Mto45fhh50C8IKAcqFaxdSR2DNZOuJYbV+lWdKoh8rVwpa8BWMLivau+M
XKNq5L4NazJXomA8td4W+ChtVfOWQVxnK9P9dTz8XpyBrDMs1ZDHZUjKetqSldki
cztWmK8+pQw0ZST9SCR9mdFnxXNgmXJfnUDD1tL2OYcelDIYsCIuwvazkWwIlos2
Gj+uk4h0h6b39QVdJiKktmsaJMyRPETVqiecoN+94F/ZQOhtQ2jaF/YHxAEoIMBp
QKjGSrz1pOJOOLOzTceKE7MLCtn60jeojQTdduZO+hhPI6oNvI6MWnh4rT+e7XkZ
AzISEkDS1ewks8Xp/0K+k7TD0LTr3+WjM3RIUKHZwzbov9nSADDGbLtaBkuP7G81
PrWBPqYr5wkFI6kOo8GHZHIsaMlDIskwbP8Uo6MJ5mbin1iAuFElnF5AYJ83Tmbz
O4weg0OrTjm30wOw4RfTIB2PPHJfCJLzxv3YUFjKFRQ3/JvPV8+te2kYTuqu7S4w
d34LBCddF2ESdLf/YHpzxiLS8YDXZWZCQLLBFuQD1fwBoPfW74JYdl41bn3ZeF5C
ClhQTBOixQijOOGVF2ju6Wct+NF2TTfhXcaeCCTGvsxV9MrBB/2T/zTFX0sd//u5
UwNhVmTzJJXXYV+G5aM+R4C19SW5Phl6fq1uh7KHGtlwjuymXRhr7DzrJ/Rwz1Ja
ZnpdbQS6obos6AfqwmoOZ9dnQm28bdRJ6wjJtx29gfwHHInyjH/fQO+GDYdt610y
NUwWdjSJnbHuvldP3ycc73Aj4jJ46CWmaxaU36DfHU8KD4dd4zehpGYG2tn7Jr9N
bKyTQ8Ary417xprIkzct003CBxVGTC9/SlMILgz+/jxT+Z5azFOzLdLx1ci1CIcF
A9HId+YYHEI3Lvrv3v1A50xh+/2UR7dvkA7+iz50ROOfMcKPp8oTfWLMsD79wn5G
u67uxYxH1vzXRnCm991GmwZUly1i8Rn8AyzKlMP9+rKTmHg3xyGc+aANdz8l9FUN
74oJn6grwuKiyaQKJ6hEuexa9M5xGykogh6SOmfGxXLRBj9cy6Jh3rLt9/SPmPq1
TTqpuivoZk7sdtmSn62MI5O6dZScMoxlHum5B5wehQjDh6FjVoMMranpA0rR3mRq
vEa6JCJzsc+oxnH04lppn5HPOvNFJ4ny2J6aT6gs82jy8Hmh4BZJrg5pb62ekO92
hWYjgAfykuYInEFyGH+VrANGnAHYdHCyHghkuv35xYngHFBxKEaCTe9t9GMYq+g0
IXCYloW2Ebi0DvKly07DZHuhOFXLhUEPw4emhDGssbjRt7RhnONetto1aFPwH8c/
vIGgFSC4hLZ54s1d6mjh2dqPh74zcYl3gcKX/4XTkN1khyGdQwjrqVdLTsedCcif
5bRd8BbGpTxFcFDurYmNOtNG2nLMsbMS50w/2Ogg64ucOms6nqSFW85d9xWGHc4S
hIs+Xlkr0iQiMXrv6uYvGgvx86xzrvcl4nqxpunS1aDWXQ0MC3Gt9CIJAywEYZ7O
JS7ai34XWW8iagKOUHI/Nt3nj0R+CN01FyRWT/lTtDUW7lgHZMnAGtELIGU99gAl
nDsTrtAUSz6km6QwDwhxfHI2hG3xOTinAB/uFqON4QwFBm2CH2PT/jZzRawArJ5n
ElV6Lyxt51+UU0n7aR1cvWp97FYDqlW8sw+ysdNyj90mF09fRhTcrIhDek0oQ9I0
QshjxEQpnUTgCnl4iY3Zj4a8ftBPuaaytz2hshiyaP3LmZlwob0L7lA80q7OUizg
7ZvQdKrkQlxqCeQCOcCkjVYD3UG3dt4RIHHInYgM/Jkp9bh0WEqMxj67hBreAZI3
d0EtNO5Ip3xbQ+/gBhTbRRDRkFQE09kGaZ/u5X3tA6wcox46dC1AaXR9//mGqtHV
v3GTG2lNV6Eghjt/E7Oi/yC5hZBQyLDCaAH7uI5FW49scDTPrQeVn1DvbE5uxGvc
Ur/RS1xjX8enj3XRke58QauBHo2L7wOioQoji5uQXHJ8DUM4XLU5MK+POCS7R6SU
PLLvYiK74KBWFymmpE4Hf0eWQvfD8t5WXA+knfy5RXN2/JpcoWrjM3T/RjikUv/y
RhqMdbW89rIV3ADs82xy4taGpAW6wYjjJgNL0BAoBSEEnHvH72z/xi7vBxO2+rLm
O1hHUw6Ma37DsjFiwjytJPZS0AjPavDcTPINBc6D4HPzMtvWNGUDC6e1JwPwHZUI
vY9aIvtDKdyhHCeU3GNpbmx+Y+CON+AunqbDkKjxzAausYasudhcfukAr3Ota67T
NU5AbcyL84UXtHFywRHNtqR3jKtleQWEF+oxghJ0tf6/3uRnz407noHzOSr35UKv
sNuHk3+9hTurPFrbo124z1h18oOZWiIUjQ3tX1ENx55zjToKUw0vI1pLcO5mg/3u
vEaoPsjgpJ1W5RHEy9wZ9HzPyDAJIZDqos2oizyI3gPOG2zCxN3IDr0bKwtB7KaW
nTqmjYSLDkbBb2bj51xkUaNRX2mNVJ1+vk5OBvofGcKSe23yNQIfMJJUY/IKsksS
l2MFTDHypvf14LD78uHDyAgla8D+cejxO/H11+D9neUXB44kk+BuYEn9Tx3uKlhs
NfqoRHgEy5cXXe8WsYSkjNByAqA7nsChAovo1DweraRKwtOYQOPeAqyc2PTm87TK
cN5OcigqWdQa2LaWkmWmxF88VHrmd9wzwjko+GFb8nsvcmEOnYnZpdIzQ2rxwz1U
c9d1VZkrSS43G9wZNtaL/CE0iquT+vRLHgNVNNRnQklreh6suSRHunEBdr8QWi07
pgZsw7t9Hw2qC9Gyhhy08g1q2r2FUB3Y66zDmjGdwrDjUg/PLCfyRReTBAOhEJbV
i1c5GU2+9xnuV9ZgBJ11N9TY4C2JGwOlabhPy0iFneZ22i5YlkvxTWa+iu+AesOS
ouIt3ial4N+7Nlzy1EKfIVoktTJPVgAzMASKiAGH4n1cEA5DlecgJsFyTj62EF4q
vCKsfhLdUT+vbso4De8bYN74zy/emSmI3dFtMiY4OKHCTBTpZDre9VhXqHrJBIAe
gigptVyNghuxonbzWAPbPbaftwOtwhznzNgs9NnO516EpD38tCORxHwhqY3dcSWK
/1lxyNpZLoPHgEt12DBQyXUYwDqC5jC1Pq5OFlec/f4EbxKUgdbimvV1wF75gLKz
TO5yXaYssPFD2NoRNwYyQ6DnFzytFret8n1qN+gU78XLwg+rUJ9beeT12DNPOKfU
VGcCFZWGTZcsW1CYKP8hkOkVJHDRqJzw+pwiW2xtJEqzGJMC/he140jRH5AyWaie
gqEqP9YdXWzmk8eLHnosvO7+ZXhRAwjywKOsv+UfbkVefl9SebwUPBL0Mzuks+k0
CbquIom9GW1nlxvql1F8qTZuLqDo+mPynAgSZf0TZ9v1DCvDCMg1aLtptPrASpKN
XloK+x0/eULfv6XXIjFCJI1/Mlaap2SmyfbJMyn+c2OIenskNcCJ7YFGxQWslcb3
UxNHXKU+O3Oer3huRNn845BPQnxoirONWdJtYIryJgdpVrDBr/ebw6P1ioxb6x7d
iE3svZDtGmX55fV8AXgjTZOI5FQ8NrvPRyvRQ8OEW+8o8abkJVWDFZQP1gmIcNjN
fsbHSg+INVgN+NQOzHehEYOIjELkxr5TKyxAIZhI3APieaHPdkNXT5sfTrBhwvUR
cenhFbOh9YVYWKdEWfiqyhz0VGGhdlFL2wwE+EaZ3gvuV/srzA61TSnBcPk1UDkW
TqXsFAtRIRVF5GuxfPveXh4sQzfubSY/VQUiop+/2XKptcXck4uWpxFmPs7qD3UH
w8NLlOIHU4jUuU++zUchUjTTkTkqoZwj7T1sVsx0bENUOQujZMh8Zz6FUKLWaceq
kYeBMVadre/XHJ9isrIiQALkDSEZjvubavdTQrFASLq241L8dGj1DC4oQWduDT/B
zZk7t+Jgh+MTo7RqPZMi6wK3tUth5gI3o37xGSKHg+sDI7L+rrdFAqUKdyGukfIn
s75OsF3AFEg8GQS8Y/2awkJbCHobzEn2/TYh+q2UpZhUV1NFFz/iEzgpNmeTpom7
XvIOq2IsCEuw/c2cCcCVE2YD4bhY80UFjW5sVbOoh+kKYk7JWTsX3uoG3hyoWxkG
R3oRiQp/BP2Y16Zr+vAbrrCjuwl1/B6PQLZvErZqFwXKRRgl38KYqeVwyU5r/81j
dVdUryAJpQdgYQe8MTSNVQEjb0Uc/rzpnjpJsEknGTYLSffsDUgecQQnGesMBxK2
yMzQNwhZZn9SxQYoN+2JfZ6ci/yDBWlj2pQYl9FHHNzxubBY918vPTcQpcWTAnas
eTCjkC3t/lasCUnUdrcayOr9gzqAx+9SNrYpc3MVnV3CRgmC7J1WqDTcVcbcSF8p
VoQFmMbtVOpswQkfhoOqfcPGhTQf9V3hUQsr6Lqzz1N9YR7D9ed6XwswCvD9CbTI
ATw1/f5edMH4j7ZvXLtI0TC8KbdZt1eb3ijrJGOs1roYNghTX/ptBZzIZmwojndV
QNPq/OZ+q8RlCnpNmLm16nTU14xUwBmHJi3H6HGIseG0H7lMDJt7G97630oAVfPP
7VgeDwX2OODfZOxiGgbLDrGDgI/ex8MQr1psbnBIoyAgfed4L03mY+R3nLsmlpn1
S5IBgD0G+rtWpKgpruW0JBvx31PVEbAr4G3KKzPPJUDxGbU3cpzEF+4XKuNTY4IV
vOr0hHZqlNVOUBjGxOJcRByUzgbOgYnNqFDYfKkYDlN+cJRLeZXMBZEDOYqvlLPx
pZoeehjyiMsP9YsA7mHywCnYMnSYVIzBqQDsH+SqwRW/iKBOnmXgi9aMTo42OUd/
8RK5Qk9RTzFREW+jv9hmGZnAfpfQ1geoqWnaJjm3d3UjH3PII8y4cdD6c7vMced7
NFCrCpiKN1GALnuGkIYR+pRjca286fjub3bSMcWXRx20jCaquA/ztMdk0k16usX5
waTLm+abEE7i96b3fF6gi8kS8INdm8v3jptBSe0E7kpi8HQAT+vooVBAs1adYh/o
/6R3rvhhfn/NIA/B+b5pdJDJqCHMSRWNp0DCeGnAitBJ1Bi2BKmGXPuVuus40oe5
woU+ItwQ22iL2C9vKKzS1qpr3ivMTumd+a7csWKu5ymfEQRve2rQ4ZIKRqc4jW93
OZRQbl9ZA6XAUpU2uLWgWP9JvXLu/6/gce7p0QLAiJyu28cWmviD66iC9rS7YS6d
YHj2M9ZMd75fT+No1MlcvxXNdawUvgDO6xFI69bE6+5MSMzHQrPy3CZH5IYuzcgg
UV5JyFzI8Ts1bHPKIYn3olQ6zB6D3efaUosP254DLHThQEXCx0h58vJ7crDGfnNj
+RuOQ/W9+7gLrUOITtuXDN5T4snu6phi9YA+exHw8RlHjemPlGeMRInZXqASTcU+
64MMd36Nh1AfmBQqH8MDIy4xqzk5iS42XucXmmBKjPCZXdursuJdXVGna9JG/85G
rjJGQaOeOC/bgLyEjUm8ms2BdX96yVfOkCmcAzXmMqhYcwreoJWLZ43rZW8/3TKI
HgHd0zo4TmeZ4O/JNjAQPcgJO7QnSKWD4u/JxMArUadWfbAY7/R7vU2Rotig8FoC
DWKU5rv3V3LTsqJKXoO6NV39gmyG3Yx3A0GF32W/S9AmUK32+Oeku8mO4b+KUmvB
1MeXXAjm3xmbPV3hV0wwJJg7uTqtDNVh3TQ9JtNVpVKh477lxc1jyYaTSGrtRHmV
GfuvhEn7T22BrSuqLcPSMhl+IewLG+AkucBUBsPcdeUqjY2W4i54KF0aYlRyaKIB
FqCxrc12qtUtE26LTVImdhL+rasgSM8Jk5gaPOFVq8YtajG48Jmh93E4M/31O2jR
eyK3iS78TEu/AJvSkQ6mIQLAcZkd8hxNvl94zwG3aeWtoG1ibrNXNLvYcDm34H0M
HLnLtAHtrnGVPab8EnkNK39xjR5G6nVnf7HS8+N7ebI5tvK09y7s0E9pi0myTiyC
QJt0t7MIvLnevcZXbjiVkGKUj8wQehsH4/QND7YgSoJiR8BYUkR2by1J2eudxbFo
Lu7VBR7KZEVyeRuDjZn7X7i6ICnrXWj3o8BHwsKG98ctT3OXMdWZ+gWD0a7G5zPr
II9zqJywr4YKSIhNou2XJMMhU48bQRBfYxFwYa5DmDyjeNhdTsIAD21jpTgbhtyg
oTAi4jZOaozQ8eVX/4xabwkwADw+YKO9vGhKNEVWUhEkxZ8RkNgVaiBLP3uUb720
pNh0zqNEOzEn6cooABAmzuPh2+DzgN4vBHhmgsyLOpkN/M0oqo17vvBYrz10y6PX
XYX40LgskqnRJFdSC3oPDbECbDmkWqr2HENy+gc27Z5yvuZ8iAKQlWDum7FdmF7H
rLVAPV/nSy2AY6bGT077NuK6S9Ffh8rgsT0+g0oBFI+2noVaD45YSUMtf8Gwr3/U
Ya9bkCcSU+yAjT6PqEfAVxZUeSvIO5bfJCnBvLuIdonpEYxE6ut5LQp4z0GeEKu7
yPTTUTyODahgAVLj5T8Q4E+BFMTso1oBXIN3C1PClan7kkVAHdO0uj6PlmENVSBs
Kr5qt+ehRqF7PZ1Shmx6mnMNwWps6aj8TyogfwaIXWmHKI5TUv9Hc1F1dr8OJfdb
fV7FLS8+w4F8gVe6tD4gqIHBw+A+4tHgWOHJOpUjOVSoPWXdZ/d09nZhb9Ug60Qe
t0IDC7bdUTO7TrK9JsrCU1C+jT84xb0FfLW841WRUbGLnKDK2kpOMmn1vYZjFgmT
PpaUWwddrBAQ+s6QcrP73oTOVg4IRvf2ZIJEyCLaBfOf/igdAWG+q/+9NRSixpkc
FuLIG0B30bSMjKXJ02feHqLyhlOlzvj5eV9IWeABAQp/K8s84oTvC+UeoCtxpXGG
BIq58Rth2YBkhQOm55PUq6cgO8iBZ7UYMAVvsdkvL1vuVUQDkS3XfUWOUXTbFCRP
1Rv7SDA/uDoGMJxfrjUTTa+jBZ+4B5hEGvxxHh+a7SUfj67ctid19AKr4udxO8cU
R1npMz+1gczNkdWnHHPPqvhKaL/3zy6YQK0COlLfwAAGpZ5oJSAICjkqxH8VzKlE
VPNhrwPbIbjUqixfRi/rXMvNIBXmkt6X8U1K0xG0HCO9Odq56K1PgUx/triwB/ph
URv0z2DTJw8YvR7VxAIBfxZOULYjIFwd7MCFHPIThykx5gYmlWz24xMjqgGUM7X3
Rim6sJ6YlBPUfcC/DDrHt03HcUGlEkrckwzhbTclqrhe+3dmnnHKuixg1SkrXDAM
fYM+wxXOuxKUF48NArQpHTHIyt/SGi/++GZxiE9U8YLjnBQ2CsUT425U3nfv5MXd
frP8I/01+wLogHdcvSWHsFByozFwraMKrHOXcaX8kApXDKQgrulXhqpIl5PUkD1Z
HmpxweYIFuUznfD7gEw2/va0onUL6Vh50ie6H84+Nz36kqvgG9/m+IsSWsZVUEhc
pGBhUXL2nkxDxP56v/DVz1I1cu8C5jFHl1mV8wyv4GmT1EUQnHNrl8P7wyR9nDUw
ztOtoCKHoBS5z2tFj+8UQ06DfQuA7JSkLjc0Kv0eJqYKlPHIHXh4bSlaADg0k6R1
rcsNDiwtCbT7LFqflIG6OHTEqLn8jFItK8dwJnoRl/Lz9uSX0nH8g4FnrSK8XExY
etqJbopI5y9CzZ0oZVlK5KKndjkhBOsIUjRZnG9Tm22ud5jRuSq0nQz65NmdrqUs
n6yzimdp4H1pPwJzHRxCl0aMK7443kAqdR2MyUpdSWmgnzweOcR0MmXAyp4dnud8
bruGQ09wVYZHQJD7b8+d1Gds/Gv/or6LAQ0U8SyMfmJNVnpVV92qOESjjEa0NU/P
m+M47y4GblrGu0HLXy/Stth7txensNcBG/f35O8tq4bo3fh94Da+njFGcNduRB2e
YHkh5eYh603Z+vAcByxmYC4wDUv94tqVLvspklXN0QcPo4s0R4IfuS9rcmI3ia+W
4vsY7p4spBNABfLM/LNQWh+owr99PthTECFqUQ4lMuUcn6n5tJlOE8N7Bju27CA4
Rxfw+Zc9sK79pjrw9kaYrv9TfuobdeQs+8/IugBLNQNG9YJ+dWrC+4HN/ox7CJ4j
uRH9x+KhF/NZMGhgnFK10FJ6FzRlI5tw9fu7ScUk0dOpH1exxsR3bhmGAhZ9fjWB
gEpvy4MxLWnl5owb3b4DZhlvzIoFkbH9dZaibfQZLZBdpC4amzcXNNU0CDMJnsP7
B3I68ZK1/HaSIgFyPBMCjplyi0XxOl1Vv77SPxNBrYmiqKpxlNDQn9XjRZwbm9MM
sKpHOUpG+qNE42oB7D+EtJMWc/DVzNpbkfoIhbIe3luGpR4/VOlTeSvxJGyH4FuI
IfPOPdMca3gcDyPYYqAvpxE0nLglD6NebETXv1v5vNGhr/Wpn0Q+UN4HlxpNvW7r
DFuEALaZYPFTKy0l9nVjYSE7j2vAsNbU/LnLNBw5uaIuqAiCFJIf1ZRw1XXfess9
EH9MYaWDAtnYAIxoTqkEptfreZLrgHZ30+80jaOggtqpJY9b7UPpbHjHeFQHOyRo
DsCEsxj57giI99QhTjwkoMkMRLZsI082RUgGzZdxde3CxwJROjIMiMuNSp50sbKn
dYqcDtsSgtv9evHXmRMSsjyIHqqmhC+FtlZ7/kpQqYn8X22rp3mlaSx1bwu12dnv
xQhwsEGBzepLNnJb7mVYPvF/ECiGmvLr776q6oZAUu3d0/eElC37JjDDceBDJq8K
N/YEDXsZ9WjTAFXJ9y5wsMUXo83aAHRAzQYPFK2XNMVWd5qd2reTh60Jx+pBscFX
12a0qfyyWZxxVxVEOpRcsTRP9gdYcpoGQP+W5XkgS3o5YhBYKmHJcy8NDFqdtRUs
dIlrGmGbZhdw2LwJRbTseymYFn5FLMJ5GfE7NLkOeGh0RGdOtOCMtuZzj8iCrK1D
iWiiMuC56qwDTWMylOC9D2Cu6BAu45OqHlsAXh4EQmYUx2/epgvcMTgRKe0kvFl+
/R4izgjwpV6F/ybLTx9pSVKA0GAuEgBGdiHOTIxOxcjMvFGxJ0VwyAx+EjDp5FAf
m4/xxoTK7Ere0c6iq/xYZNV3kEYV6eOKZ+pVlbTzEChbLXFKtDYKXkfZ56M7EBSi
nRsBBMvz2zHsqlwMcAy9Hu0Ds0rTpSiluvzZ9xbX6W7vQpbKPSWqNRrnZdpPpf6g
MCHYhBc2zwK/X7zTMfdxLH9IgjHw7nKKx8KaRqrNwZl79P/lHCiqrl1FarmvAEtn
W7eZPjlvMR3Tb2BVjFZp7EQOBArNBM/KVtD7eNeZktWYm6cFHmhZ+flsr83BB4H2
rU6wk086ztKsczeqeVQt0lJa7tvHnB7RO/GTHUig0PzHPqgeHJykuUMI9jaS3uIq
m/EoeSpy6q4AGdp3TAQ5vf3z1VAENdQXZfz3LnUWzIekT112ZDqVbB5OO2otGJ6/
jlN2ANMf1jM++sj7Lajr8OsjVOw/ckzxQpsk89EnEknLzps3E1unXMkQVmjf7Stx
sTg4wVuBrtwVMIE9Yh32nKXdRR1/tPOq0O+CLpLINb/Tljoj5ptD7UrVWz5rE8oq
aDvj1PluTRUagiju8JEoZD6ORV6IDAGX68CZmNqbOQrM1izLIqDF1oYQNsnU0UYn
3h7hI4scE5ntqbzDkpBvlDikVpFuOoTWmoOr7b7ulD4q5bGtYirS0SiF4S+93PaK
V623Nhd2AoI60/2GtDLrwhM8/WBbXo8RwtnzRkHjf0VIEtGjGVbsuEpuL/W6WTMX
CyM+zm1FyfM+hwWzb329y/2qFw8SDWJ2eq5OyUQkh0UR/ShmEftvZkHD1p/FBfJx
vwoE3PtlN+ZYiKuYue32uMBpBIEmgW9ynSTVkGB+Ky1xBDLR8ZIGlhyl12foCTTh
o6TyRgLaWVa8HWliW9fII1CLsbOgHZ5ElnZGzHxDJvmfyjAj1GQ2tS/hpeHnLTVq
1PJjH6H/4ULUKpwXilE/8bO3FsmXbsPyPRZAqF5bb2ldSRl+ZROn3DC7TZdXaBAT
RuAbrKtwsBL32ErjsHFRsuMCELFOeMdtKwhgbCTt5g36afbbeYVuTidOqEudG4SF
gl4jkRcICh1BGnEiAcYFRC8dJuQprz2EpmeYiK2akyQpryM19Prn2zSx2YBlfh89
npZIwam9T0PAAuT8Odz/VX/poAgMhClKorSCMAAHsJ8w0Fwu8MEo3qpkItcU/awx
n+ubfyjHArSgJRhICgZwrb/9DgS1iWul9f5TN1rFQCAUYdtm9H9oMMu3PvezfmmX
/0+oDucPd3AfmQBrJdYGDvYPlz51SVIRqVDPhoLGogrFhB6aa/CQeOZS1pQlTr57
uGrkLNOK7Qyv/z1Ycx6aojCQonj6Cj4wF6Fr76eNuSeA9eeRRiUxMjy8Xd4RgH8K
s9H7ZYDz74LYGjiKgtOLpz45FbZxTZx+5HwMS/eFtNGMWTXz81kTAJYnyB8XB+tG
Z8jziAav4D/XcOe6cvQ+ozPv1LwkBUxn5t/FAW5f3kVb1e4XON4wKOkIYM5IGRHH
6tV4Ai+Uz1h4KcygwbpvCXY/NkKcohulntgw65xIkR9pq+yXe/FxfLSUyVAFH8az
tRFnlZA2Pfio9BUON0SktS0unqCImOZIHHlxIWBgmFMmsOVQaytc4Jk9EI/NBq4Z
m7XubuFYFlcwr+ktVFCsq3RPztffDRQ+sLv2Y9ERfTZFn0amQ5vzS2k6gGxrVccj
ldcsYBkLoA+EvjfM0WArBOHDcDHGzG2lyX8d3EHo2IIaQzv/sTFRv5gpLAuEQpQd
XSr8moYJAtQIm2l+cPbHHY8q9C9btwPFp/5FXWNN6VKkT7asI3HXnzd5Vkc4a6nr
F+fC08kTt2BFzqDe/J8eKp+1DVUq26WGJuMM2snuWYteXjHLjRySAm61u1MaBiAj
vAXN2YDPWxOHHIdfvJ36dW5K7LMM2vFDcYp9UJSwuda3ySwB2rgd5RsLX4gz1lWh
aXDVRF5r7MdecanW4JaNwAGJbi/mrCJwEI5lQx2/gP/airoGBL2pnzIrvbx0vL1E
xzObeY4BtcpbeHYuj0okxRV+jGyJ8QIJvvtFmlgOaZGGI0eF99ynytVSBAU+2tSE
LBo1OvlvaZQr3PB05pMc2rkJ+u6oL1XDEoFElqYAJHf2ZZyW38eCh0/jPMlhuT6b
RswyEtRijs41Mgzi2GQFSeinVpGTMtDtqle6TK+8i/dWo48F/LFTOvb2HhzVbv9t
BzkEbXHpVWY14/6/+FsdMHbUgXKYbr4uE3Hu5Ervza6xvgMGT2WAAEbo+Ghfvenj
yVrklZROU/weWZwBq1uW7kIVeNKi/sUpHDDN7DPz7k4n67lsQ9tjdFVVG6r+LxQN
/3HvGxh5p/+6RikV7U330wj9Zm8Djwpu70RyQdRiKtRoTtC+NAqns4y7zdznufO6
0hIONZD+r3T+nWwANyoHYKtavjKrT/nly7IWGHDio/2Dii81r1Gja49dLSiZ4I8K
T+DaldRfJH9zB0nLcemB54gLTA9Fb4fqPislZfaNcXc/0N7jTGKSq9zenZUmDA5+
rJgQBHmUTFe4GlrI10TjTeBRiQSiSzIZbN2x1vNRp2DhoguPJeKs91pQ8pHJ+FBn
b36ADKFfItz1MHJXxliLG9v/GeZryEJnXS94F+nICrGMRt273fYtgej+8iZ3BQm0
KWKx0IvIhe4SwmyzEKx2s+mkHyP4XWglaNYHO1roKBtpLGKgCfeN15aejhGNMn0/
WBjnYVEluBbt23/dV0hHGOuYobcQVexldhfeVcU7K4wXQ71j9filfhHC2pRt3AEZ
wGxIq6hcuzVhxkFQ3t0Fr69VOiqss6fSyOUzZcp1WQBVDrmbkmZDm3bkmNDAap1P
g0hGU1Td8XlJaXpFK66Vse8lCY8nMx251x6gCZAE/PHlAtpzVezmjqITw00+uvsl
M9Zy//3poT0Ki/OrOjQMPRbEaMG1zhu3w4A6kmydeWce6lXxmA6jZi9sUUaPNpd3
d6kDf8SgeP0IRLwD9CGCRWwX74XCROTqMuv27DXC4m52KO5UcsMFZW7rH7U6DY1R
hmyQAMIepFDC/WBMKrxx0HFkaeAZF/DwF9K5XZ8tWFIsbPJ2wa4J/wJujOmLZWPS
UJDYoDzm/Uin7D6C+0XRlr6+S7C0oouv7PjG2rpLLTWcNXwXa4ktEEFwXttjPdUc
GvLf0G+07KubCRqg7XW5kqrCAEvxgAyHLK1oTi53x9wUEqu9G8+c6y/KQVkOM0iw
SgznSFN3QdP62HVdRX54On5WnxNHazMvuZ35BZTMPytk8FiQq6SQyFMepWkl7iBO
gTe30NRAOTUbg/C/eDFaSzvnhqb7nX4a7qs8dK2l1tnwGdrvoE9ijgXSgOsnLZhh
vUiSWGINqijaBq9cyAxTNU6tJXqDJNE+/Ta5hm5rwhEOHfAgok2UXtdsl0flZgi/
m3XZIikY2jkJPb16qjVB7IZDJkn91d2Qzlz172lhT51+Qv1o4g4GdPpgtaPv+fqm
DcWaLvLOPk4CJ46+Vp7M7B3ngIOUp0Unt2nd2y8CSbXXzzJTDkCa3OAXHicgNXB0
Z2CVFipQKzMLO0S/YusT6GW63wZM5uXSJSoEcFUWIDZo36wGgXfUrckO3ysEcK7D
Twh0lbWTBlpkTpyUEZ3f8dgBzlF+Onp+rjHso3xuyIVEQXd0c9eVJ9qOTMjVYrMB
hFKKz2js9heCNmALqKViwzgnFuvoOqEtK7gBZsfMR4PRgcBTdYnQHHFmpzLLow/L
mloZVp5YaZvsNwqn43S+jpn6IzPoVWgplEDbiCQsBgsmw9ct589hFPYZHFAIYyy3
wKFaZ5vF5102yH68WYG1dc7fMW+UH2f0U2ir9MJoEPytkRkdZBcPQJUNcfkTbEUG
QsbveYS/2LtBZxin4ZKUfGXWoaDGc6nyV/bwOChl71gTE2uPjYzWwbKRSf0VhoH2
fcNXo1hfrCYaKW9fPNYJ3QxcHElbyJ6WuyAlFYRoU9FrvmELCPiG+oynTqC0rVLf
1lXaU6owg6CT3uU1g3mxj5dNRriATamkByFlTRExW8A8QVLUxiLEx2QkAgfyIU1w
eJBNZ/nmGfA7FHTEjmhAXS1OSeOgiOlmN8VDpxRcgeo46C0hd1v0LwszBUkub5w/
0ZbK+HIzxQzEP4RfIDzqYYOasm2Yc65uVK6nO/PJlWqbTpFMg+C77yLozS3Ln/em
RskOUh7B+B7McA+QOlSAHXh0s+uuaAi+wVBVNF1Pi114RFY33P+2q1a21yhRPL1D
Kpow5yvBWYlagFrm9gco10HUm8lKXMHpzpY++rTtqHY2PWtqzc1RABVidK+/cyqM
3hMLtQPDqwYpNUB1oad8kPmqPuO2gZN6YIgLLMIOWfEaN42UCBEfPRCtsQPcVWoC
RBozvpay4vitbyDY7Ul0uxs3y4Qo/FOS9wLXvWlIM4u95F7HEvcsX/82QrjiW5YB
0W4QtVLAlz7UyuXi3V0K2Zd3asMmKdhocwJBsehN7+3Zx8HfZd/gqxMxA/MjonO5
OD7uOoQKlwyjGWL9P4igQTQRHYp5Kz5sgghl/k3/eRr/bUgFRkpDjaEIY8KBlbz9
19vL7XSm1Y2OsG5U9FBJIkFmu7p8IdR2uJmLnMC7jRSeeJssEvfrbv2aC4Gr/bsE
GLl+nZ/ENQ2/Cn1JLDgIMHRDEwOUyCMhDk+pgRdi2VNHepJAM375xrfV1jNiFu16
hoUmxaz1h/L72HqQk9OvOGaFUFlP5hLqWdD1y1sLU7lGT2OEDWxO7G4StgOR2VZv
+HCbaU8qr1L8nO6wANfTRzqPnXaV+B5kiEsLq7gDYXfX3HcfFAJOukU2qNJcQZFo
I54now8iU5gm7GyN8bFDBkWDjadwEbjeAuDuD9Xgsl+7fZmtJVco4VJmeE23UInR
GtjmffoOpcBAh8FLuQYEwX2zuA1HG1uiSOPYLdQQnYVr7lDq1usySYDEPFjpHhCh
d6ar0Mdw+h90eTJs1qfJneKbeNWNu2j31MDzsa8HeYMDE7BDRUGrVSLPbj7uOMnF
TtG+JHnJ9swJm21TGarpxWVIQSAHAR5/2r+s+kVf22AEvkutgekgDKCQXfy0NvpD
OX8N/0E9IseBDg9ou6yOMYru6Y1vU9ZsoRm9v8QE0HNtrdaxMcAcQhX40d4wWFNn
4e7V3ZjU2xid/OqPhXe+PQCUk0WhCVvABs0Jokr5u8hGA9T0WRv73AXdt7T/HKrB
x/K6Et63v9/1ksBqHXrypnN7blTMH8P1sXYv+2MzDxXeBJQ6d4i8A1sTBZ7LtkJC
ZGI1FgTkWZzTJCuqzc414pUyHLh8/pS0ukTv0485H0gj99yYKPg8+PfrWsqXT9RE
9b7K4STt4RHpbATQQO1I9rWHshFfZLMf7my91iRVg2GerEwJLX7PGgT00e6AXnOR
gTJ6dTOcO6er2uvzkUkfUCu2rM4FH83wM7X9a5tIlNwG9kT4BtqZ8Ls4ouYTOYTW
oBfsfO/mD6d7NjeFtZQdp7SgnKpxePwmJRpS0YmvOZ7P6naOTzptvGDL0VNPlYW0
ZX2r87zwO1Ck5JN99gHxDqKDH+Q8aH63peIH8+qys5x+5TofhsTArp08dhrbabdW
/Qru6LEdPUCLuav7xJG5XU7rKrt//U9f8rButUSMg6rB8U3jV1bhwYE9Bp6mD22D
PD0dYcTOxo/0EuyGe/npArcQnnbc7WM0igRE9H2X+qtKmW/JOvKdwguz7lCTPaZg
Fjkvws5LY851NlNAaAKsOgYT3ToTfatmzRPD/6K8mz0nXDcWodakn2KJ1fO3NM5Z
NKyFi4m1wAbnxeJ9Uwn2xgYTHk5NWRVdHUADEWH+x1EzOW2n/btySWyl4IbU1w2o
XUHYsIvmryf5EovjRtA2/ZvPSLLmcBUB7rSJKFl/lt7dFFAZx1fe4Tz370xZnPEN
31bvcChXmdKQzkXoWNZG19t0k0gvy5yVWAeS6GBhTck8uMMFpWJhNuDS+DQhds18
twQsFKnn6l2hsEWLm1vu3G+uzBm+6HAVAvMKuEbtNRalmLZMXqzsLSHw39ZHT6By
93VnWtTRkRgN3yC2U3n8+obG88UJLOR37Kpva0zk4XkwC4zxMREZKT7PStnuYVZP
wT3rqoiyQcRThuPU6mBD6WeQKxmOOxh9hXm383coz6hhgTZ549Smi92G35fbs/OM
cqm3SnnKczXAJrJO6bNv/qgGp9czft+3whETKda0QfezeeELgpJx/rgFZD2YwRz8
NRuqe9EMrhKTj4HNZP/Ktl7zYSa9aCKv4rGmdWsD+SqALEXKPpaR4eH2aD34j4r9
skjWD8hMalotgDraqp3DWFzFmCi9PazsYkjoPLVvZhK9qTdnyq+HnGaMXT36wOH2
gmv+VgNk+eacz2kx73sJLgVRlP428VXMQ6+gns7MKsskAxi3uHHmxBqHinB8/YAj
bRjrwwx3bO3x+sv2l+cZ8BReG7kTP9tgBwuqnPHq5xirHuSeSppMcctDeXUI4XBk
wZPdBd5XDrky6knsKZoHoTLLtYmWubNldNTQcj0iNbeSFfg4z6hxxxi7XkPeWgnR
kfEcm+GAjetzJQJz1parNggDLG5vR8hpH/KxBN+GhMZOJSQrsGP77jfQO5IpkH5i
8AaVBWF76poCpaUSd2uzvAYw4JBUxZkfx45M1WTHE4PEjusqZ+nwau37/3OlzwUH
yEnfsANqG+DUo+CWe3rG+XhcOOOoFzIQ+oANb+28pxJzwq1Wg2Ym9DdHX4CbHt6G
Tv0QfntKPSyNddbMBzebTm9AFwZlz7CL/UX5Oz15qIuFMTScdw6q8vAc29fwicbP
1LTtTa3nf8vMWx6uNVB//Tpgc2REfp3e9oBdCVnbJ1uuIuEfWa6WU6QWNiFbQDRx
86ByFmlthSSvIUlDP7khoRzSYAAJwkWgIhKKNqG09/KXTxKNNe35VB2fJ0jDE/n0
5sNkKRANe3gKgsFBLOwrADZ5Ntz7+bdkdp5LhMnLHxlXp5igDrT/XWgMZ1kJ/Azr
ldXjXD11u7EmKvkV2f6S5N72n76LF4rDTXLxd2+r0/PLV4k4BNyQBTXbDJ1BHqQX
2Emwwh5prBnW/A8VaGa/rGdPAWvySS70MNwtxCNbrbdLMQ4KwTw1gaOBWdAOsrIf
8z62JCoI0WK5eUtqTRuoOJinrPsVFzjKhDKhpMYUB+jWquGzGmId/oHnbLwrKF76
BwOjbB7Q25rQ0TOEODiknKzCGziwksyTy5vAkvL7PEpsQ6u/6M+fPBnhX3CPOIKz
0Ve3hg/S1EiPbD/04sChrQWgou2kX+fmnM0zeHDumDiaQ9fdXQsYAUoEyokK0YFO
xZ30m1RKfHhiTihuz771LuiM+NqcANyAnSv+EtF2uv4vq2kLPTqr6YjBw4aWpveD
3eG7djixG4fcW4TdPcbDDtvuXy3db5eiO8Uc0FY6NGSHSdBfNMJD7LYk2gPXO9ra
cXnnT1u4QXrVFClpI/yr7w0Zgfnzi2j2/ghX+42bq/uSg2nPSDpPFN4nhVd+8XGy
kC8AYfs5bUBnATDvDi8JPjZQT+HVeNtHkt3FzWAKt0QweX5BWdIv0rtriweHZLOG
bl5cFOsnrZdLqiKH+cyYl2Dprcvzx95rB89nmNERaQnRDezNc/SolPp6sS5Tmdt2
s8T9RIUw4lq5DI9B58CR8aoXwAf8DcxJYvd0UxKxAKNrCF4krvYqFUM3rxFz0iSR
0jBamwm3UWnlnWjqjnOgMAT8t7jMKuEiJIAHm/dGIBpsaD67vd2yAVBBGt9KqRm3
L4ILj8U3yqn6IhKOgP6kHAyGoUBbzYM64eda8rvlF0xjAXifmzh6BVp7Nb/bc1FL
EFCfbqWOKDHwS3JGFp56OF0dHnsXrAT9N6zvTgL4BRh5If1Mkd9OYkgCkmqD8GWV
YSpq7qz2UaIbJx8ojc9P0L1RqhyrhF+15WwLea5AC4JczTrJY5DfhLw+6VAnrZkt
X+yOTD5ARcGA24pfv9w+5AwXmUOizXOV9MAkzn4B8hLPbUskHYH6TRaPW4SkBEzD
NdpkutRXhgsGY8KqwtpowSNL+vz/c8vSN/A86IyExIfFbeAXbA2mucvWGJ4M4ANp
HJH8qUUkkQBMBg6A4AmlC1z83LmX3H2zr22urbt187mVYg9gIjZE0R0ewZor7Mut
haHY5qzbeRufUvMijW1PMoPV01/e4BeptdHer5YTcoOBwymkpIGdVDcyxAy+bfU+
89O11UDkrMO/LfGMsrmwvqZfIsLRP/g5aAD9VnTsQ9RGQNEk9jAJ4XcqwA9zDuH3
3Ajm9w15QJDystshlkbQlfrIjZahf6dUNs0zfXfjZKCCcsPsB8e3mhPnLzBrNn8Y
8g4FMil/n0JY1d8HrJAhpKgYEOFHGS5Kr/iuSstcAis1m5bASwLxbLYFfCJ76peO
2T52IrLPwPSgZdYqhFaRpYVVET4MMTg68KgnwencPkk0xki31HstQRrH/Ea21Dwa
+G4kG/c15wXsYPbPn255obUllC1oKdA4iaf6+hryehRNgHJxbeDNLLU3wZQ+l3fD
qu2LfbTfmoctH6elouBDCPRnYRcIJ1DIYbJijpuZs+W1MjnHllX3pUHJIRlW1OmW
UMd/VEHJ4UYGi9IYRobfwebjX3ueWTV+AL8k+ta4KzuSsyjAvyEZgT/+0k9Ddlqi
VKgJcap5pRptmF98kefetJE0BZAXNc4j/cxw5MZa2iBNtjHSEvL0Shj5lN9VGhHL
wCBFjGZwRqoyWyE5cS+pXiN7Tk1D3rcuRIdKaKegJsYBXruSHfQNXn7IuU4dzZJ3
UUGsEHhaqwp1gZGE5X+JqIqv3T3XzXmRMVGccMRD/E721o/lU35DqppxT8Usw3zu
OBMmu+WPVDMXQ49Xu3cnCIBXuXCBgImwj7PSslLD3V3GF4uOZ5AQDLQVvj4XfIvp
7rgNS3jC8YUW9NRkviB2V0sdOhYOpDdqmBH43R9ozV4j1JUzx02BESl+wsMal9tI
4jFCgGCrA2HOzIn6GFrgkRPco3WDT9EcRQE6nXVlPciJVMSilKVKDrIUCEp0QzxB
PrAzgEVRdVqoovGq3KnN6wmV7ze0rnZ4VRcbDB1QbCzCqbYa9eW/ZnzhqicCJY41
vHNitEnilvdpvKFUd5x2fxC3nNBsudwKeJi1gZTI5j57iZWe2mO65JHeXuslDk0o
kxQFs8dLtITpLs8cNfAwqSfnEw0s6FhMzrVK1ij5NVyXydDRlyzhLqC4VN4LOP6l
3xxatZ/B3vfdQKG8/bZ3nmQlNZSfebPVhr3lYzPPyscurj5GXGjNjfXAlYW8bETG
oCGRjqqhjQdp9WH+KQRN2ndNTMnAUqpQ7tYOHn0UcdkK//o+7qWKRYg6aoAbZkbH
zKJVwc7ped7oja41j0o80garp01JyujdQpU74b0rX+PXUXw3t0bCw7KF/2TyIo81
mdPr/Erdwi3XuVqOpPgQWuC4kn/I+47S+XtHRcjTV6AtwpN9h29NH+kw/nQ8rQqi
expln1JU6Xw7M7516x3jklYDwsehHDRYWdZv1bMALJr1QJHsn/GTdzUMgG40JINu
5ZPL9mlWDGUXpQOx0KzrItUhvYw5qqw7bdOLPUAhldOtTahb6kV5aNRekIRnpqQf
cWqqOXrww+LG7ImjZlKZ0YoYjta9j+eaeU9SsvcgOeqTPGPE/OFReGwzHQFGR0pL
6Nqex0iUaY98roAWV9fRMvp2iU5s21PcO89uwTwlg/XJAORTuBhvEyafFcWPbhDj
RcKsCH5EgNk9TiMfRCawPBhibVWdce/JgtxtqvH+R9R1Q6goOqtxiNiyqnUFaLlz
HzfZ4ec7qAOHmpnqQOochqnLSYILiNnCLHRPancvRQivRa9avTqBQSr1J8YvC/0f
EIs+vwAuGEzrp/55C7l15M9w4ZlKsJOzojCIt3gSB2p2lzVbKG7C1JHMZ4ctZ+Oi
/V+csbhzfUAUnUnLYCBRgDLlSLX8eKfecLwUGBd1ABlcd2DTwQQJvL/iMtJTims6
TsNeZJsEeojFPu6YgdJuQsFqgQIVRvwfQejyzlAEs6PlehKvsLJipzR3Cscipd7C
Ump8q0MmNL5qMdy/eg99qypWhsFP3pAiYDg2R2r84LCoEz1qrxq2gllu9c6XJP2Y
bE6q5lCtcmsbNG3m8g8RIXXQ0h1R1o5+0UFUkiobvtFWDBIlKqCScvHJaqgtRkxm
R//KZtArkQrBHTQJ06ixPE48YuvQthuKzGgsCl1uvcbkHmZxok6BqQObARYgOdJf
OFzCibP/x/qxs1ifO56jG8PGfajp3/BosMMv+fr/7Z40KRnegHcWUNefbypmF0Sk
LvN6cO8v6kastw5YBKwtlZReyZkRAqm0fMCI3yAlrDGRK0nGh2N+hk7rjh2jwneV
brFzSMFbLwtsJMMStyNZj/Cbr7Ry4n5QN1aAal4MUbsqkE0ZudjhZhA4Lxf7BsQ+
vyfh1GNJDcZ5QrD3inIrDmLK7lTH0L9hHbkeOBB4jcaO2s48PEkBG/7lLyTPgbZz
Ewjl+MF5rYS6ld/prXS47Y3Tz5KLpbGAPHNWXj3mitpAAmhfPOd2XsN5BDUBjrZn
HbNt4jfmYZg0XtdSAwOKkpZplAxFEy6M3b3sg5WwAD2Q2zacljVsLOYKt7qPqSFA
MHugaxNcomgakG3fM68Rs8FUEoEaW3f5sPcPksvCmwPNiiS4C86ytb4I4heb6lLK
GPG5zKC8tbVtFRiV0hXEAqpFKO9cDslo/0PB1f/dInFvldQni13rAnWJ0TPbwqhW
nEiq0sjkOWuYXij0xFaSalrZ0Yaa9qWWZD4eF/Wktwv5KyvhIpGPh8cIudNCYP4I
FoenUsdwv2k207SqdNs/MH1PAWCHBLMPPUB3Cr60rq30ey2lgj/9DTVE9j4NOoFy
Ii8nayIMT5KAC27TRAV8nxupDyUwYGIGZmwkHgLhaXC6DxE7DItTbtht6QyS/mf4
AT+NeRcHkQmvkAaehGaLuL5tIzzepaQXBe/tMISV/eK8asRJpEIH/Yi+4dSVq/2O
TWHx+sIcQ3ZEk8rOH0MNlu2DCj30Q+w6AXlmtZrU4xCfpyRI1D9Q+gtciMSiWd7u
qpclt2XCUvep36TB4h9jQTfBvQrwyd1NJHM9BIiFwzJ/JhZ0i8GRM+nyzABDgfIZ
KZRklyegdVJED7yJIYoGa12x2f35/1lcMb5MuJJ61oQWH4u0UZSkP2aJ1nJQkZEy
CdMaciz0rb2kh549LRRpjzMqr0Yk8s2eKhMgHVDSl9jvETclM0LMmeT+TxX+ondo
UjNWrHIdIZJRe3jRKVmqJR4laMm/uSiSlSsDh1xiTZbFfrkj7e4QNigTXpQJFpHX
rTDM9/u9YnFPLZKqUxrQrV9gQQ+8ccv8VhvFWKvSa2HKuVHrkK0EyJD6JSKVLdab
gy477aWGYk4VdRXq3EiEkHBvS3LtV6j2mZGLvyqZ+oxeW1guTI9nWVyHMgX9IklB
vgug2w7J1WiXr6pXpfWIoFo3YRAIMbJu0yfUsljcQT/BK1MFv59xYNp9qxYXh7dX
jW9i68GvPHeSGRIPNyGiMZFHNRNMKtYBA7ZKu+acVwgAF2bak4HL0DGNKtj00O8s
RREsiWQMdcfdwuQasUIOt+Njx74G/d6BxzxChcZUuJfAcsHj0NOi0iRbcjiqVRWs
YIsrqAaNJldsvtgFPTw62KKfcbhnUsQ9UUDp/B7FoGfx//f+gUgT7iKl+3xZxKYG
fslWjDroPvuiHtlnoULIpPIO5H3u6x8FnqBspNchRJM2MGbpkHILuf13eSiZv6Ca
e0TqRhw5FWZxxVSsmzFyWaG3m3AThXn8uY2Jo9Pzh31lwFSRzLKUu2yKFj8pmNdn
rXeQwFMXXJLqlMshMiKu+UYBCLjOECNbhkdBz3U2juJRoAY9y2MGKkQCO7nSlbSC
8E8urlXwKHK4wowxThZ0CMIDsBbJWOW8Uy/NaAtoTKhQW/8Bf1zEgUgjk/T1w2eI
3S3Tt00n1jhPi2cPLn63G8BWBsvxrmd3Qq+ozkS9M4Lcjy2ODozMFfj92vI++UFC
qUHAHs8PR+y66RilK8gVYUaCDgh4ovYBqjUeedXuFqbWoOrY+vLB4MdR/BX7+Tjy
lbb46n9dJ75SXUXvEl2HNbhHrMf08TAPU3Vhx7F6tX3crHTDOdS1PKeAOI1TWYd8
G/feCf5px8jEnk7qKueNkeNZdCS/DHwDHBM8CKO115+0zFfGjYXQiAiRDzkX+o5U
PdT6UobmPhuSZV94vKNxaJ+VNrVtM3Xm9nHxt+GS7vyY+nGWXY8GfQh9/+OB8S13
sIGDcNfU2nM59F5wCLEznHqiQaNPv8ReeXTZX7pWchqZVgPwIolgX8g6+9cOo813
woEXn8D6AgRk24/Lpc8+j1Upm2MEk/FNDfZvoQrTxqXHU2/pO0WMp/LsJUH+r0L7
xSDV+WAfQgrHXT0XBr7dRDKL+O9KVEazAFN7MMHXRYWjJuyglXXLunGABPdXqM9f
beO2K+m03kX7ZWL5HYAUdB/uHSbyKEaZ0z2ZzyW3vwfzSx4QoIitN0TK+FJWhMhY
YAUohsLOymZ5SnSrR5ytCRRrvY0yIunsNQyB1Zi4kjodavQcAEqJg82452Xc8hhn
a4uHXl1+HoGY4N6ZgmvD2pX6XME9iw7aD1qCPNCVCh/jGSDItH5Ss9UyfTDozIBJ
fmmy/zWA9oAR4IHZ8UT9XR2+DI6rQBDMaXUvs3vWOhiUedG9f2DN5MNn27KoDXe8
0g6MKFMco7Nhd/kIaKe4yFGMW4QHD3Ju1Hf8qTFT1nFBkK/k+QsdADGL+GyhOrWC
w2MUpu8r/SBSPevEw3bqc1WrhBXCL9kGHldsCayfVuq3AOZVWzw7xLJqQ0gQo21v
dvSVCxk1SRfbv/Dni/U7q4/z6U4BXwfftqowSKZ3d/x4iFO//+351ebp4g5d7d0F
rTB1DWS5QMrotGyCyYika5Rz2Qgb/hwqTD74XKXw/qJ1goJjx5P4gNg+AHkRSodr
ZKMk+2p60mpWk14bqw9u9czprqOXrdobKw4K7T0YnsGUXZxuJtzj1HSwtjOCqKr4
R2j7dNKON9SfObrparxiDiF/41CkksH95hKduHxDsV+X9CmxGehN+gvo7dtgIuLe
XU0ReHaEk7waTS6hmyRQ8s9t4pUlfUBr+pX9hrL40J41rO5xZhvTkMtRrBcmUrkG
8X9H4uPSbWHJzOgL51n3IL93x0DfgwVlyFqPBymAbKrPob3GAprmdKCwjdQ24Lpl
qowBzJ59fYs5Ob/UYyHkb4TJsESUs3/A/Y3x3Tw+RBa7Y+JOhT5RKtcoZrIolyQI
cHUUHaCwDWeJp+JvpxSgqH4tdC2Y1PYFJk1eGlaf2BC6/AhyEu/2PgE09lX3VwXE
sSBFq/PKQelr8bjvm2MjOl3F2p4o7haznyXd/4E2wXn+f2MUGWRnc82GJ5d9fnM6
gJodh0XjwrE38iWHVl+Qhl37OybqPkR494nTo5LzYeYY6YV9i8dXoEt+nwIerYlA
WBVRR9vlK01fXJkemUUIMdIOJoTP2UtF27LtzB7ty4jm3Fb04Zwbx/0Q6EiZFKvB
kL1GAcV7/2dQLYj2ygKJq1c0+N7fwAyZTdUDK5MLCCY8/60EfA9LIwMFTcR4Ptx9
8+lOXcc5OY4yrWskRoVaao+sZeRLN6NOMrXMbuMgSaYUIu0LyMdMrGOxFtYwkT+A
DEb84J+sB2+BRwoiqx3pahl5Hl4i9clOW837XGV30zFgM5BoaHbkevenEtI+kama
LsdvXwL0nRyAwf7GUqrjwoMoYNiQl6aSH1NopnoCy/hLmPkOftngTqutvOkt+J6t
wAj3HfDDanXUAiDj1nJbjEH4/YPetad4cLEgfqBNEi2PYeHbR5wW8CRWvT+14MBX
4Afp2Ofu5NOTETdvii/mOiD7Y9wBYRBES4fVnqcvJgaMYdQHHt573EKT1iopwsDl
NvbZhifutuimpvs4/ARzSWMaXyZTEw4XmxA0b4BM9fRJrG8ioi+1meT9Puh6LxZy
oGgyrSebhKGbujNwpluDDylsSaObtv+BhDfn92rZL30siZ4vkdwkUYv3vus5T5+w
889f3c7s8P9U2G4VHsT/PmETFutxbFo0sfGSjzX49g7ABik4UYkuj0xNGkM7/KTK
CA3RlB3Q3/o2VXC70xZnc8R7GvVW3wvItMUEGDRNQKV4fIHe3QGImf9OfW/hbTso
n+jP5wZ1n1Z65DCLmprOQuB95Uc85IwEA41FlkSJKAazdrBWj2OV7+BKegRwHykZ
xSTlFFOdEyo2GT3r2L076FVMhBFabuSVznIdycLYKm5unV/pUmcR7R3qiqfS0YLT
T+ZT9hfDi2kWCnZXJMMJOR3DxhV+2sHJkrVZ5l9uFPyGsMCCxwuOl9UKeIgKSWac
j5hclAqiRpL2VWV3Iy+DikZiD0Y3k3GHIlfODdoEwh8S4kpuUDnBZPhXCJCV3DXJ
OS6GOcblRnulJeS5HdnfdX+Etg9bsc6gnhprRcMYC5wTCwXlZ1J9t3/O5K5nGBeJ
42pZAfB349bSNs3ijZtzpjhh97UAvI5Fk5mjuhfBiuo16IASCeqzQgHf1Fq4zRiJ
t+st2vsdvvEYrLhaakHOwGEpAvSm/dWv9yxEuWTQ2xNW/bt6Miut224gdhl81rP8
3yk2M+9ad7Odzh/jqAtBCJyDtCN8vq+Pst50Zj0PGah34AchIe5jaySqlpDVBOHL
USVq3Y9xaCMSVpVJyMpYT5uvk8asjRFlKV9iw2cLrT2B+Yt6+vN3jpILrc1PovyE
9Ds92jwtPb5/9IozeOi1y22W2lbcFFL3N1J39BxZ+fq9RRgtd5tyIhuNfL+n6fRP
VRO7M6rzNDCkQ+jdWI0tlMptgDNwQonXU64+eYqJ9GXs9ofnkzpDk4tz9IdCNJWL
bUpH7bWqcW1tmdbFrqiy/BT3vvF9d4wbeSWG4m8l9bAuOOvCUY7LK/drt1Db9vMm
I5RCG25SZkIt/MJXIEieyPtxBXollrFLvyXAZmNZ0OmGGX4K5/jLcRVqhvpOPh1j
UNpIzbwIWTRLAYtfHQigTVkbgIIIa+O7hEZRUDllF9TiPl5H25i12LC6YxrSwR7t
sHF5BuhfkT3Lqfgrk2S4g63ZdHhqHh6DlY557MXpaqnvblDJ7m66+vEVcG+B9H+A
E/tX4rkQLIMgoMTLxmVNepHX7afP5bIU7T2gYs93A6l4Sw8J1LS8Nu32PRSrCxLh
y+hAIldfQtBUCgVInchbnk0MhnwLA8wmXlLS4htYpne5W+7XT5XWD/QDqTpwTv6/
uAtZqe9bZZzOxx8HSALnb1VPJsRANhEtIfk/FrEjpnPqjW+xs12XEddhzR2b+eJT
8paTcY4sEA/hBqpV0KYJe1vpkV726omVJa7aBlSQ0MNDLI/YDU6MlpgPlr3aTeUH
BfcAMfeh+VxpC0Z3FjPG5WE8G+jDG0eI+ARPIvTZagOTrxolkrJYQOp+HF3x3ePf
MPrVqmzw/CO2910azlQ9jC4kmesYtaVpOh/+l525NKF02cePVx2unv5Oc2Qo+AuM
5L5bLeWkt452A47f8hgAj87OXRwpd1UmUoLgAQlvfSIlHXGaHy14MWKmYqdeE7FF
/AgvfUDZofJm6biWGcA6xrYcPJbkqdAhVsyeN3tXT7vy+fHe13Dx/WQ/cFnWtzu4
/VD8fpQtTXuPf6fqsWLzjP4MQbBarvWvodoBACf0RdGdytfoFvX4DHlTdVnJYHkF
4r2TkXQBBIJysMrwfAsqc4jdIgwZV/ywKcCH5OyMpVBEEdnUUvWTjmwuZul5O9/t
F/0ZdzMoUyLO7ollINwfwjHozITJ2X58Q6QJiT+AKLXl3oifNJ7cxeM6VE33rDZg
9ZdbCn/l31Mh19t6FCRvm1ZknQlom4oy9QSo5fW9gCr/Zea9IBAmSDf8PLKDxmfD
CcmZG+y6Blk6BXpC3YHwEgRi2pf7Lip0Wlus8otrnSt4ug6oAa0GFW2sLarKchnP
3vAvIYKJqegx3fNColsdBkrElLFHGQ3Z8KI7R0cyVr5smn51xXlOXzloaVxetZbC
gYBZ7dgsKP4xUYB0Z9bfMPe7+hoqfPhW4pLh63CO/f30bjTGPphMNUpVyjgzolB6
cUynBOj5MfflAl/apJbIks4mVCnWKVzbTuMUouX+OYiPbEtcDSP6L44DeTKdP0Tx
jIMEg0QnR/XGUuR7uow/4csEr+dEylLbNfmrhi6t/PT/qUo/SRSiuhGnh5NzzLqs
z9y2C2yeEyq4q16mJVqnn7t+ThplWt++SsG20Qz5V2elX2cySiEJHo/jtBH6FTUk
6UcZZDlWm2vtCu28kRnQnNJSbmgcCq3yaeTn5Y03YQrRnzEBkO4zgRD4erxoFKyK
oblK77W/XQUh+EQzHeFM+4gxpGWVs1ju7deadxmS3i89gQOCkwTUMQToV/R5z3wV
cu7KqiyzxgPoDsfR/wQnvGA3dhhb7fX20FlI+o8TUrN4+gUkGCIh/CWxtusJP3gx
kGppPm/MlGg/iCK7ViEx7u9TIwZ4Wop8Pqnl7WJFI7+v/5IcbX98MqQSfnolQbF2
jGv7tCy/CS6U8gb3G3pW99N+Z2XSyTJLYqkxfBr0XCDsi3RCStgP9hVrGkE7HZwd
MNGgwFTxfJ0t/c536RZ+qH0qicwnqORpqIESVqINVVBwHDlCyruwABUsyW9tPzEb
9g7nZ9XXwhxrYf3a3c7RrouS6Mmh0007CWwXxArRgdQJHs+ZIVtl6qeoeZR7t4QT
lCFf43ADEiVlzLGhgalwVb6eKGytACf6kqGdB2K2L1ha/9bZiIaHVqvpbA+FOHZ/
ZeEo6zgH9CeorKK+3eV51bCRWpvZxzhve0Fgxc5XCdhOkuEz+RTq74O9feO4uF3f
T6kJ55jEYLSIanwzMqw9ymB+l06dz8R2hpT21btSXsdAC1IviurDzb2vZpeWOj1k
0G3fRMNXVTnrOTZz7ihtbOROVPBaP8K1gPvNglFcFOMvkfSl8w3Z0PgMgG25/Wc9
IPg7+UDvv0O/uoUZNEn4/4sagLQ4d/sy/zO6XejRB667+rk7yZcoAsUaWlxqWI+Y
db7nVEKBR7oniwTgizDjWKJ0u5t3iii96doLNKVbcLaLKIEjiya7vLUUhHYoIugm
yogXwbuGUpxH2nFV+Ib7vP4g6/LUdBKuYEp/LbSxizglsSVy4jaVzn9wpuNKXZBW
Y8phRVUFbw/SuDW5/mmR3VALsnVYVlKqLWggRk/dif3xk2ou8E0ZaLUjt32Sc6Z2
JKGsnpqOAR1ZUZgRO0E9hfURm8OiUMRJJmoOB+ZGk4LQrBs5rkGZ6JW0ust6YLN1
oHJvOx1njyej1D8zWP6dwpzq68sZ/2QnBxU3gdCY23cdi/C2t6U8cqhGuEA4ZTK8
JrzDCK2MzJdMKtAdDONEg9ZoChP2mbA6yB9yEtglb6PnwcwlAxjHkq+E6pZKAJAj
4atKHGUsDhzcFptq7NtR8Ri1CzCl8zTCwxgoVKYvYuqtB11clSalNJHh0J1RJhd9
3ZyXI6dSnG+LArqlS330KrTQld6jfrN3Y2X+mNqGVHrEXllHigjC1hS0STeAYOEi
Dv4HMCNdcG7TBzHV+OGoBoZuEeZJztQJQaNptEZx66dKrE55tTvDBGKoVOYGAEw2
Ab3oGlr3ELl9KB10LoWdwgEgtHLt5o6P7tpf4sHlrEVm4wfQsKlwzwDPVR5+3Xv8
Cn4FlULfT634atWdMZXArU+AkadgospfPEDpBZH/mWimdlvYZ/eQ5doqk/dduXh3
Vj3SrvMuLxSd0YYHIHPF82veCVvJgUnHGsJqj1CR7wP70n2Lrw3xt5+kTD3XgoCd
PKdpaFrVxtPFEQcOhY4KenKVBEzD09kDjDZw2jUt+jCGOaTxswF+L8cF0yODJPKZ
ePzdqbgLGf3qweDj8I+ukxg/P9QQIf5M2zAxspXBY3gNucZjZ4yS+JVibShdIIR9
M7/kPVZubwlv/+T0Rq+S/qdH5JNwtMCNBDWh/iZmvYYn5MT+8UEqQ8yfc6b+NTmd
AdqJ10GS6xgYGtZYIAarlnO0Kk3F64IhX/j8bHt62pGEoXfRXMJMTQaf3NWwcpAO
Q+kzm4pdc7J5Eik2PU7afl1x/H4KgcX+CjmOrGo2XGCfa/bdlNlsItSojfa4yOll
nMU/PwBSWb2IuH/05Ojy/Wc0EvhGBaHfzEqQMd8gTDdec/ZK0u74HDAKgQzXhFGO
05sBt2f8cPBp8uDDJco5HPOglKOD7OX4+9Pro/Jdy8O8quZm0T4z1T+oB0tkQfTD
UXTncYHOVMWMyGzU3TM3BpJKtKG6PfAS/CmsxCYisRtIQO7b3JtP5R7jaOYMmFex
5Pd6PnyvMmzLSw059N/NTJGfRAoQaMBF+VZ+En7iqynRMJHaO0nholopFNRmLU+d
l3Z52UvQAGNMO+bnrlUHtbfWwnEhCcGrHgECwjTGfDba2wu7X1IvTI4f6XvazRS/
RRNKIo09/w/mYmHWx5lXecRbGNirCbRskTDhLygvHWdlLvK99kBG8vIKUWUB6xkm
1tQ0ysOhgp04I7QorJcOBf7WK2Lk6m5DW0yiRWtFFA0JXgvVVrDhPUHiuCPN9U3Z
+dmlUkaVuHFDiXltVzyrtQQfgeVAkhupm3NRXffBP+tkJOIxkayIj+mWm9iO4xgG
pbZ9RJCKiqGwACNe8kBCsk+IYO21ZhhOLStfM0xs2UWe12GlffcclFFEfN02m3di
OSiRa+gdJFWSQCxIuSix7raC2VF1fU3ISsZEKpJmANnPks9sgB3LAcENxuE4k2Hw
li4ltvjcBYBFaKiNq9j7HJ/6Di3iDivktBl38G5njelt+KNuYEJtHiFbuRNkce1l
jEhuF/0QAl4uO0F+aNhyMfJg92AkEZifqQBEoIBGVvar+qfe+72OTOD1/2N2b6Ew
ud3w8q+LczQ5HbIcPTt8xsKxkSVG7e3JCmFD/R1UXXF30YFe6jDfLqGPQm0GK+sM
Gk7U9rdYDoQzgT2G5sMqS0FFlam0VbBmJfdGzcOLZUc+yUuh9upw4zGwDHBJYfZd
9Qkn0tWeyqm3N46YZZb8bhJnDR37ZUmFg2oTmn75E4BGxAR3mtMybDxYG0N320wo
iB+clYB+cHhxJ4DbcvpwMpAR6YdNd1zmjfH8e+YiPlB3Llanz2gnLQbXQRAV+9cV
lpjmI3t/1mb/xGHcc/nia/tiJpAhS3+7aTl93uA/uWTldJDKltzh467XKHZ/6qOJ
NBPtPwBEmrzFfhv4vSj/MZs3zwk7AY0EdiQEAmpfXLHzsW4kDGkn9xmJi4iymxKF
8sii4ocNXKNGdEdhF2u92Kc3KeRn3bkmaZdG9tmPYJzFhZHoikSRu5+hcSsIrJyb
DK4g7+wr2VfN1yufmZldE2376k3lJvyMCNgSSUAddF22iM2cxqpGShg59impVBYi
1xgrw5ExJncFI4Mkcrk/sUZt7G5Che0YPMXiU+x1JNkpbzLAzGe/icN7feXe4Ncg
h7p+oKwMUng8oakwPFjWEcuXV1Cw1ZNAbAY5RaUsIvcT+IzE9FqzAoXxqZu/tG6/
GGQu8RpV4SgE7WAGlX2DjaaKTRJVRp6rhUpxWAngT5FfG+0InIuml0v0m/uSnBxZ
7T4/GL0UMWXwCM5iwhJABocH50mt0R1z2m60jc+hvM965TtSJxXmZsk36z4LR6Cc
WYs3EDFAOLoBQTfZsY0dcbZn6Ryl5KONrhrXh/J4odI57atj3YPoF6xLhqBDYQWr
wFcsEMnSsuQZELinYfxPURvI2bReYjQqC/Pjl2QEkei7Vadd63Z/8lUJkLkuat7X
+oNChwSCW7TV74ZLRrqPHT/ukzLSAuo3TGE7+DQsXKOzIGCSXHH+9YcG7HEBJ71e
Z/eVNO/OcqsNFe98D6kYNd5pjugh5JivZgQthyZasL5JZgXu/2WLNZPZktQLORWc
XWxNzX4NkkeI3wyxHn3xKvB7jgMJheQbQhYptRC+yYTDkxyHE16owOSPF2k3HFD0
59mxNm7o2NlhQiX+yoFM9QKWIzydYcludYYPg4spbJHMH64q5vYbdmKyXCajFTTo
lWO1jVqWC47n+OdRpa6ao75qyN6zXQgbWFgOUke0L3qbwTW2LgmiTZ1nA3eg7OT+
IDe0LHeSUZ8+odvEcKe4/VA17G/qJ4SZGoD+GHzhSHjWbrxW6kpJmgZTkgEb8ozW
XTxuDil4yJ++MXayydTrfy199pci+yl3uDgC+y3zlQr816gg4/v2CvUv8hG+vuRn
0ULRMrSNgyVICttSbHzLjjIGk11p3qyWiygua3poTRLYYmhGKiw19EWrjc/F0vrE
XCeCQzp1iTB+ndwHQ3nHS5traU4GCXtRwBgQrf55LsH+KaaaWqDAstM/Zx5W3pqM
WSpKF6GkHVbf1VBCeCh2Vb0FU/6GcG3EFUyy0UR+PiOGScqIH1ql7exES7+P8909
g7pbhpUwMRQ3zqVoXcTtES3gEBn1m07bk9ZZ6zIx6WOeMU7Q3aurENOgMn7vZUMU
E0LcwrfGzHTPdXxFqDABf1a8aN7Yln14T8BFIn81kncte0KUPKS/8RuSRVYMpOid
KWKJDRUhTUXfuqCP3Q7n012y8xxKAUy9hIPPncj6ENUsuGRjAiZQyIHedNceMTLZ
q3IBVJ/RcyXTE+6Dj9/YFEFoLa/sOO8rf7ZMbYHubTbdasb1c52n3Xr1JUKZnhkK
sfMjf8ablEf9nruah4yPFD3Ee/Tn/2oMUZyDGID5/nPI+xcvGm78CpOqmM/QfGZn
ik54dNF4UKt8uDl+NARxpEvCpqGxW3GfsAZhEA/laBG/1W7qnYHLVkajGA8Ldg1w
n1IJU3uBpTZxEvlDntL61HriIbxx31wN3P8rZdUclQSx/2eK85jQH6PKYVPDlYcz
uSPNhX5NODzPKQvL0fyPp3eMSE2O/QK+CFxhPNvbpGgO6E+JbFnuDUwDPq9uJsmo
9YoRDheMnqxNl6ydIanQEGVR29D9N8ffGtqyW6pZviMgOwXB1WXKataOk5sR4tkd
sO2eje8SvxeGp21tDB711PB8pklcJga5F099rFPD74NK7T60qIfZ3P5DDgzk0//0
NuhRnLvo0fUrjPRWIQB8QmmD7s7TNrjEUXCHlENhx5PM82hNIcjN3ZuSKb+rGvp7
qImpXAesC5BqSVR3ufrCdfn+H5ofgxD9n4o1Tekc90ujwQv5ZcUkdb6oa9YWT8aE
2E3v8iKLucXvU9B+OpZv42OBJkUwpBkpvJLqVvOSAfNqpLDoIHknid+Q36gZAHKd
zluDfn/hyLIsW25RA85e4vJ0eyFCNAQBpGLsyYdAVNd03SVLjfydUQ4gyVZ9M0oA
j8DQr1stvKYh/hjj2usDfQd1gv4M19QX0AL8SPXQF6fHKofAe3/lBIz0XWkIGKcb
CLzd4VFUSeqZatTtnSANFK4G2dZK8RiHXyEdwkN1gGSiq2LPaomUrf2q9FBt4mVe
Joui3uSO9Oeb1bxaLynoQSTTzQ62LAbLlWDltRhiUzwMtgW1vs8CHnPCLg9DOUI4
q5liwn/CB8mYu0vl/W6nE3R/7fOjLVTnTDHHT/Hv0rOrq82fRHCq25rE+RG8PZc2
Fuvi9S8haqyCMIh8rbsrPIrNjYOIgEYesjiwfAOvqbLHEVPMsN5WtTVvgKq3k39c
nsbh9Gj1rg262xATK+H1Z1B6UOpm1Ah+nSxUOW21gwpBY4kOMWLmTpxLGaF9j6YS
hk3Og7vZeljPKEfiwHrwQ1DMKYUDhBx8x3dMeOsCBKyJr2BehGdutwMWHyH4H6VG
UqzXnZiAWADwj7a3Q+ECWLeEmPRYTJU5SV5iMfmqAs2U8FrGeu7GFSkXouvNhPhZ
WmXGrFKeGcO5unjd5rS6aJs8kS1teSuNUlGzNj/Oynblr3wUCDMv6bNtbQPMnetu
fR8ilid9X5MUyNYWUeRStkOUj0LVPGpORcM1l0Qie0bYtvPwHZG3E5zy0el6AbUb
k9oOXI+d19KjSf0YwXgPfZA76arkjkgtN3W39MV9haRXsgAyQ5CaAd739BbMJC7v
PhuxJbihQUTA1mIDvwgITRQgytCLwnNcAv0aSvJqX56ohNcwwPhWtE5s2Rx9N3tD
JQeZwtWXiBrQrC9e+W0jbIpgBlRw+RvnSfrGTHW7xoYlxX55PxwZW/Wjfx86n5s8
K7NLg5EGe7uA66lq3Kf6iGgTTuMRBLLwMOrGU2QqcyLIyjKbNr75qLLeXMUka9TH
k30UKvrmQwOnxssQvNaLPLB1nP7fC57d23mhAVvrrCA5VFIPnrAkjgkhDDILe4O6
ffra4q8rrqwDet3203HKQy4slbcKwge9/zDqZEqgHEv9t8mVJNf1SQoLEl0DjHjJ
gCXF0yBBGHn6STvE14BZgXVLpbtLV4eN0NyNFwhad4aQ4aU3P+NgEaQu+XUziFIU
HO3wwVSCWjuCM14sPlymNYf9BoJ00Vs0BolT95lzKaCdSC8jvBsczvgUSdmUerGt
DeydbP9ubUTAj6k4OXbn4M75lDiRpoziIcDuKv4wEwXvqDfhzkPkviTCm/Cf3ys4
K8RC0KxpO5DRtNlPSmW2zur+8wr9DuXo0X1WkMPDA0pXOM7pLGLDyK2GDPqjmv3q
IgHcvfZwCrUJX1AL6qTdz/1a8Wtk9pkycMubEwEofRzkGWpk8N+by6AumyEraEsz
9CMmHoE8rGPxx+2XjhdQVTedINJ81okjE/IW8nD5NLUf+sHpHscBrDekq+5167wo
1HldPl2VkETh72hIR2xf+4ycQW+SX1K8+Brn6nJgcvrteWi3z9D2X8vLXprJfjmg
qXmsKXyC2ONdnsqSH3rems3UEJ2OqActK/u1vlYHoD5bv56UoP6TkD4MfpZUhogj
QIzBeO0+twzk0EUT4I14W+DvrpJGdDUVF8nIsW1c9t6d/0wSfaIj45eMAORtq8R7
Mk7a7jVuMYjXuRw1oNF/UAYjpj1R8mCgcdeOvsIZj/d1r+MiAKUgI1BOTbAQHSRn
xr2rkfPVAUT1A2OmPNtYzn9J1WjDCGjYi98GnAIOpO0xwnS+Tu5yB8ChASWalEnr
vD2rGbpibBu0ZH4LtvpuVGceUlZcme9USxlKpXWb/wdhWsCUw+FJNftdLli5IsET
Fm5S8BTzSTfXK0NqfJpri8ysraRUrSZQV/6fKSmOpaxR8Xlt1/LdTgKhfDMQs881
0CD2vPE7rHaW06InvR5DryJEeQTX+Ws8tDOK4y6icuCaXyLu2Ss6Uybunn1VLBYj
Ai7zS5bcHdp62XbSMINepq6rcay/OMO5GnKb1fXiMlSviwWXRIc4cPoMjMZOrgzl
iXKsKkllITuLXQ3BKLDhm6Dll+DyD6sMx+LSWp3rYZKtbxgX/wbuhHsS6ypAdV9Z
+XEGvFhk8Cm9lrAeEMpCCdUbFPMAHY2cbILe5ggo7LrUS5zT/a4fih16Uq9xs1kD
mRYDlc9agLsYj577fEVXnlIQx5ExbQByAeOsUAkn9H9Rnq8hpNCzU3GqEqhVed6d
YQlm+ojD2CaSuOFybKyN841T756h2QBmyPBfSDwcYUuiOtpY42nHA4kpkEH2lFqG
p75Qsfo/+9ruhFQSKu+VLmZrXAHHin96QVMVs/ca1LH0/hVSasxsfdyNkjf5e7Rx
buoKTDLDoMb40iTR6CNxoDXiLSlNklBREnb1kjpTW2Gtn/T9K4ZF2q9mczOQIHdy
baYcDc+R5vMimERcUeeY3etAr7T78IlssqoIms9x51Q1xjR3vVBjNzdhiHtE7GDZ
kuCywov95Nq60TZT2cvtPTGPVtHD7IClUaMptWKV+A2IM/h8qv7Iecicuhectnz0
72BX61dCLtwyArqRn+grR4UmCFo2+Nvm53isxjdt3YfHkJZE5We4s3pdZGxvVs7v
pRU3wgrvA3vOctQqRQT+Vx+3/V/znyCnjw0tGzwgwcE7CWcL/+oA9U0xWOOSwiUN
ENrh5dF3FiXyF02xLuf4RnI8niXd7b4cnk+sQ0a6+ePjt8GKTBJabHSuc4KUbYiO
8MpXDEHBYJtjAVJKC0PgWA1yWnFuFuKjBaLK0lleu4JgszSBsiZncShmYHmP5hjD
dx206FkodAzHQqlGFQO5DkBTEBHqTUa0mDvob0LWVFO1aGGz1ArklsRuG2596+I1
n4OwLrsEqggf8LpQYHXD94Jw14vKRKgaVn7yL1dzkXzjE5aN9xk5W+7+bQSQJ4kJ
K4EFv9YtSSEFQwML7yNsKPfn/z84R1qTTrPGOZqFbvigkjY11vMhZl8fixUXbM+6
7jZ4S1ofwQe1bkBSr8NgoUVKmjJkZ2kGTJp+8Erklzmn3QCeGSvokYB/jtCGrDnp
KNgDkYgBiU8olN6AtcgMcCijAWBUUdSxhkUDt3NPtIpP+ziKH47zj4I255pmov78
ZhNMqWZzgjPL0u0WPyVFlmIyeEYM05kx0mt8fy0c9jq17cThnnGD+1ZKKZwCE7I4
n/Y6Ef7fnhq3JuPUxiCg4qeY6l0nmt+pf2kEt+cN19j9z0bC3YrXuwPTgExZc8YN
EiMeYeyyrAaGE4t94j2ej6s+yaV3kVIGJB4H4mJ3yWPucLExRnjFp0q4n9cKBL/J
OCH3otoXL375yFKqyBkWOj8rqpbg3wzxjTUc0+GfUqKxMG91PBvZuw/afNg8VjOI
0HlVp0qhgl/KN3iKiyhL+a6BQfZ9CizPLQwbN6aa2hVvYqcwdPeLikFGqrr7hKr+
edHQYTpkisqdxCMB+xeqcgVjaL93znJUFFnZLjk+LPL2bnsRqmpR0dstDKGxmBhR
2/a0CFMLY3KrAhkpeLi3IE+XQhegVGVRSzQonKn5tN0ddqv3ZnhH6sl+u1c1AHQ+
GJO7zlAZA5PteNWsKMWlPut9zXqw9oF/M/8k/5i7rCSbZRYF9MQuCmK24AZf3lGI
pLaF60SBMzzNAKO9Zxg/iiSu5I+jG7FvgAEAPhKO5X4l/4crjOUTL5BauvVRhPw1
LSRBT32mYiYzCt7KPaI9odT3g4QAekZlk5R+hcMKsce270ne5inVGW0D5LJyN/5K
Vdr4AsN6xK0Y4CsvwNxh8IpQSpLSpvL0NhLcsUeFCrg9InMCvYxHAomExiOK+51X
ibJ4F62Rav+DAQe0c7Zq/VF22aLhvAxvnFezcj1qq+ABg2yWpZPxterFM07lqV6F
1tCAZD4km9qrZGoya9hM/uJlnMENQyeNjfztD0R2rmutXD3zGKvhHnOaR+R9XGAH
6G//BDLKekkmIbWH/u7oSWpGtm05fpLbDWKlnsDlMcxDHwKB5jU7JC7AXUSNQrSA
gTFrdzcbmWQyrxfUVlfewRZ8l1T1UYrIIbbN0tMgHU4iwPz6WW9Y9XxwnU9++9ZM
e0V9ueieE22BuhfUn7+RFgkBEkIKLkrCfiq6VWzS2YZpoSDo0jn9aao3/xZfVFr3
k4XxVaIwULP15lVAA2eG5jF1Few9JQZ5XaQhYOtO/i5lIxs0rJzNRyB80pwLMNzg
VQ1Ny4rUgVRDM4ov/49haAGHMnYuqH2hRrLxwNCd6PwwzC8uThn02H14piwhRx9W
w9nKJYdqluLl+3fL/QLtSup0Nd1lnF40IPb/Pze4vwOy3lhHNKXiXz6B3ux22e6u
ddI1ebqsie2D5B/7iMasplwcnCtujZa4p5CF4MY+Ua12iGviYsn9bC/zxWbh9oIi
Upu9SZWchdi53rLJbj2mUFDonJ02s4IBKE9Z8dOXFVZb8ec0TxHkoHT17ARpJgw/
CYSqK6Sj5CQBc0EuI5lF7qxriqcOMLpkDCrXN2x7wHmnyQ5qXQ67JJzcMD7UUnS4
Z7M4/u0A2eEBq/1loo6MKdLW4waIwo9dtO+myhxkSMyknsvtPcbsLlGR/TYLt0jV
lwWM12msLAXzVx/lu0BUO9zod3+F9Y0RhUq5tFBrk2V2pcztckRXe78V2YwZPIX+
5QQvvr97sn1jdsCyDUKfu8Z8/kSGF0VrRbuGgltvO1ZslGUr8gEGVc0OHUEWnL3j
ihIv/fikKYEsoGvsMnAM6jnrx5HQ53gekhv8+W2pYb89yGOxiuKs5o4OMOGvwkiu
Bxhg61gNMbqdk5xYmE81ByZuWHLra14EOrlxaun+eORa+vrVwGFLo+pTZXaveMXZ
0tBU1YtSqcJ/4ffRPxpBFmAJndn/XMMHiVOznsOVyM68KS8h+PQz+rFU8Cyia3qq
iYR4VVF8LywOsVO9lvw/dO7T6wcXts0prwFnYqV2fWZkaed/e9x9DTFLxDkTaH3Q
EmpeyRNu0loJi/A+JRzAtdlR62m42HUNeveL3JEgj0t9fSydTstMCy7zhrEby2gJ
fPE9TzzSmrGDjex+fxvZaTild5avw2yyfhK+ifHKBSZ7d1bk0QjpIWGCUa3DpyfT
zicBAiq29BQF+fijFIzR/NogWB5SJS7/N6KiO030jm9zzAEr0Jqzod9/Bcp2KVDr
TXGBzGaiSU7LBGHBDNkHj8NXGjWP3XNsOBmVbDDj1GNOsBehfqo3B6Bvn/cO9Fy0
HNK0VMNu8V38KuKM7r/LiJHwulPwv80+nC5IIA4NOwKvSFZDgnR+vTdENAV6IqLt
OXzIS5ONPw8RkXJB66jj8S2lPETkUVTHsa+tQ6aR4rrx9ipNQFbCZObZvbD9sPTB
Qii1OdFApKF+/J0UMoVnnhCg/9KqIo6CQR2yqOlhCv8GY9P/X5EyKiqAljakEeS8
M8fC6M07pfHPApnDWmnHugs2MmLp1kKUZPYBriywSAHzDtrJhpY2AOcP51lzAnrq
T3pnOGT3n2UU5XPWJdM7t5wsIgRldF19bTxi8otMOxzKGlNx6KzDtaOEiFTIUkU+
f2SyBbEavCNC9/jpb5S6KxvqLz3XbBJgOzci/fWRiV1KijeqX1CogA7HgERPwGbK
Mx5DeAXCNQAywvWdiX++1C5O5agP0MwcTHG3ZRTcu37CBy3I9bP/77mWRYPAbSco
ICVHFhQCSl4/980SfuxOCyxWtHPMLobQ2dv2TvbC5hs4QaLPzqeAsYq85N0fXvi2
yzBdv6HekKNI983Z3My/mCk8Oq2k1lKVQmfCbMACCoF/la+9KE5rG9ooGajwblmW
1VpznFhTSrvqgu1IfAQ/0YB8PcF/b/sLcuYGTn/KpeWQ2+SWdh2tMbCtWiOP3MBM
l7Ka5oEEYRuBXL8AUeh9GqPSy7ZB9zK1318LogYgGMbm3RzI4ByR6G3lnF6tDGwj
o9+psNBGrDShqBQWTJ/UeBitp6hUycrz9RUdlQW3ctSjl1+wOWaukX2rkoZmPvUf
IXq8EV1mdUEWSEG8ES5NgHcy2iho4SadpEJpOEf2Vp6fJUa/KBlDPv6G473HjGA8
LR2SNgFQ3nOViASRlAk0GUYpVhx69JVXJ7k+WPFXkBQGAlnZS6V2RYi+Rces2R0K
h5vXcgl1QsgmIWHOemXH3hgTxGA4PEOqy9KdNER5LQbpSq5pdiQKUeVQxOJ+tfZ8
kCh5hzaWiUwwDUbk6j/3sgrkPmBZHyhkWWfQwdXzRpuTOMW85X1401mefyRvb/Gk
H8OcM9m5t/mYeMEsQQMulCx3wDueGLuHT2WFqgGObvXmZSYLxQv7f9vBc0PkgSe5
3dR6sUXwrJUbZQD7wZWMQcfL2FopR/yE3Tpv+1HTvTOE+f9Q8EUyylnAZBrisdO0
iXu+CQOXYlr5L544LcZYqGdiL46AYo9iXIQ/NElYch9pBd8T9wdbiLVhPk9yPAMW
t3cn5GFclYhBvMnKRD5hHKYct21mFwj53zLsu+cDCUJ1IH+m3qqmAVrsuV0e32Ae
iKBLaAQnfx+NGoP8kUS/6p7bSz2fXC4KLzRixD0R7t7ZKAJ6WF+I6LK+lknM8Wtq
1UlNsufVaftmaCiOxb1l+CusX7ZhyA+B72jkJGOzhcIRWiiT1ODuFySvBRcdFC5q
ieBRZ5v9a3Wgx2DZ/e5xr1/uVbQBJRaRCQ3drNtd/MSbVKICFQSJGASLbHSWo6ai
g191dsVDZ8uJjj2rNBmOrLLUFjkLBgHVZGr1utw/x8t6IivAZyUGw0pQtdGfsfwk
argHOR79cF/wKH8JTC1rZeJWSZt/utuT2owmsRAh8ajdccYYo291IGTzLwMizBJq
ElNMe7RMVEgZtMyIzDDxxyNwKGl47E1FpLn2fUjHXrARsR6rM+A3XdYU3b3vHZUz
UL5hh7zQ9v85V7BLUVxTgZH732YHwLVRqJJwT2tJ96QyVWH2Dv0W+T1wnsrKuiI3
FXH19Q2Rw+iVJNr+pRMPmGvgSmTsWiMqZ/NWYv2uQYD0YIP0ZZkH0+GLGGYKKqlv
ZUMoukmuixDGk+fyF+bKvScTCL1BVjlLr6onhd2fNekvmeV69zaAwTUCsVNMNTDt
fPMBeYJ+6NZfxYVxVIzlCV6qPwvPYSlndTJQK2VtY+pdV8sl8f4Qnrvqri1qfwZo
SAeC2vpMyOCIfGvqOMpJUKG1ig6CFmgw71kv4zvRjLd0+9wXQRXvOu5buJcqC0dX
yI8yRL5oz4iNOU+honQTeo7RHFWJBUOe9FaAZE7oQvaeAnT8QmrhEt+hGKwI+0pf
VGG/eMBAF1wRs/xnG7L92Mw3X6539vaE6iP+z/xa/Eo0KQXgcDt4eARGuYo1rvyq
+TL3F3kKNxJ06iZryelpakw91xXVEgf9WrLfaIpZCjrxtCWz1B83BWZH/Z1IoOeR
qGIX6iXGSWsFl85f4rn3N39fnCvg35sVI/lWp4w7fkpuxJ3DpqeV540ZbW+PZVLY
tYdeksD0A2ouxJ7khRGMlpGrakh7bNktQZu6jvAbeJAbuNEAvp56sZ4PT0cDv0pK
6qOOw2q2ZkeJogktur66K8d/6lS6ZCp/F3LaPBntwozuhpk+2OretwWkkFfh99qt
Ob05+CawWub3uvXIxaZtRMXbql+Kvxhd62jban1zxUln47zq63PXxSdnXeTYJUgL
0p1cd8f0fm86f9TWMtQbulJkSRSnkg4jGgMyPlCQyEftoaT2ueJg5hDXCEZ0v1hV
mu0Hwa/qIXXoqsQ12e+Ub7muHDdZRbEbtU89QGMqB1bAVWCpxLcV3kcwYlzPY3to
0Bm0L6eduUr40pgEgyjbRR2pShzIq4+izhXJ8tDmSzAivXtKkykFyP1EvdgP4We3
mPm9h47ZHJTErbdWSN0q3sA7digyQqPiAWnk9ztGWjPMt31bVVK5gUEFLPnWKKEW
PENgYqZyey4XIllzcGMD8+IuVvt/MSpGSwN85CrgoXjWCpafF6nqLuEI/MrBiUC4
egtm/mLE788Y0ge6nLmrGRytjogOhjQtHABoAvlJiOawAz94Tcfj3cH/4H7T8WeY
Psd3JkVkvlAht9vChZMkeXIgJ7yUx0faYmDh78nIKkBbpYBehXiBK11Sj6xEDZvX
fHSgaYXh6cudK0HSC/lBYdM1MWbLTyPPLOl51gk26UEHPb8qPTfSONyDvMmCk+62
MRU6wJF+H4QBWrfeHZEptNq1hsx6xHB/LH85FKzq1jO457bth9LMnhkjE85YT1Ze
RNH2GaY0ihTLz4tma74af3wGOqQt2ZskuXxhsuh3ULtt30MECZKcy4AR9MLrESxa
/GUcnnrYt2ZP0RSg+Kaj3wJuT4xYJfQc66g2KwGJE6uu0Q6RognzSng9S+DBYrhx
+INdlkTjQzuS6x6tpnu8TeJXniEe9IP6HmCerrwTuPX+fxN+dYTboi9fzlP2PE3W
CZXIb0oICaVFetksv/v0ehmd1dBqoQQsHNxl/A0tilAv0LYeBZMHAjgT6iqYT3xj
DKCJ3IfYgr4XG/V791YHp0Fat882sraz+5QmP6pzncL3ls9OcKFckFR3xod3jhPF
trId3VrgybS+JuLUXBzoojKhORUlGCJFoc70QieV57ZL70nSJCxXElhEziA2IrKf
a4J1Gakv8NMELgWejH9PWBVdtzbkpn0G8MRaI0DVnGO3jfVQTC1QVmyjKBoRarIL
Q/dmJGAo2L4iYUW2HU+LaXzfAPP2ef59WGsWnq0qm44wEFc3Izvjh+KpcDIIRT9D
0UrvmVNkkqEe7MXaNyxqKNNU9rl3hdBQVgjIhdj1Ph4PCCA3mY8jRdiULnBmFRde
l0iemN7m+r7ZNn04bVbivffo0iRzFUyRbDXnCuvmeynf5Lf+QuQ3LrUxB4AS+C6a
PmGQ3d9OIpK/jXsautoMb4I/jtVzdqsBtchgDHoFoAIJfmQZQOKkc+QyjjXrcuw7
XGWY9dP4tqFg/JitBNomG04KDei4FTPoJIvsf9huovo8pJNcTst8Da1653x0RXF/
WtEHuNOptVKY4FSFmdvAE4xyjToD/je9KT/nQF0wo2lTC/69D8lTwA0Npd19QB41
0WUcmgvvwVSSGzDWCNcT6zlVBY4N/1EvPUQL6OnlwURcPK7XgfV3pNlsd4stEVjh
EO+dG5vFecsd3539fDFWGm5sq2iH6mggxNB6L/Kn/p90SqNUivOkNhgvYQa4O1VS
Zkur3COd1yXqjGL93rSo6Noomntb3CEv0dYdn2ztErP/Y7nElzBZJ62YBA4EtqrT
FHzwr+9eMf13p6jMON8ULu8HDihec2VNglb1ZlxryUO/vxUiLmuSwXajxWc7X0lN
8ULyTc99VKIW2CX6SyBH9ss7gBxjljydzmmUCSQaA97T8KXgz+0kFJDyI8ZB6On2
L2Vm6HNQd2ui1r6S8T+OdCwpdLwTMUbEPls1NJ2/Lm2K+yfJPoXavp44v7FvXwov
FmDvzoKcfRYf7mHwiSsqULGnvvGp4cTVqbhUwsj3MBj4Y/YOIMXDFxb7Xt8PsGjL
kYwA8Ga8mkrsTMZajFE1f3pk5mIKWF53+yV2TgpJIfoTBKG9SB3Tn7Bb9NjVHS9B
+Va8y+9jEMC36wlAoJgjWVJGClP/DuCmOyqvmODM5t6frzcreDxAhvCnjr3LerBY
nuOP2cLLBP4j2wshKvok8tecESCV/ewKmrClQ5qxxguyqNSGl0PzkJQrUViDNNSg
kyuhgLelc6O1qxGJiS0sUVQ2knkdeYa6poFl5ii0tz928GV+fx862nYxJwEGoScL
TsyBTXMCmuFMYvDOEGFwhfoSG0DCUvR6Jvq29Eqi0ePbRtmpBLZaGbgpaSsJFveL
5X9zFqGNUvOPZA8aKETqawv5nIdIMD6JOxKlcLMHlKdfDg7wPhsEAvqyJCFVrho2
5QplcU9bzKGgviUFDWf3s8bebObOgdSi/WpAclprz/5OkC2k39wpvpQHQjfPn/+l
ZufP2yfwaNpGwAj1lDQQdhizI9rS/R48GhZFH/XWXAs+JMW+c9oTkx6c4pB9309g
b8gLKQDVC8tB8Lduedk+64MqNy6sjl0eOqT4XzoqUcH2Yek41mjn7+HYA2OBXl+D
j0faZA3dVIc34LoQgl4FZglm149B8ga87AIDDj3UbiTvmcKXtSAeRjyY57S1rUCZ
ti+rGYg19GfLYaTy26e6Lhuj78N/jUKtkJvw6J9JFiQqYQyH/Pep4IA6kIzz3ceo
Df7jDuiHqaXOfPV4GH9RTX5ey2SJ6gAP0KrsiJpNVLmJn/E+Jh1P+9K1g71JZnT/
gqsdA66JvZxz47ehMovJEnpxiVVlU8DRPh2DYVwSxZXB8p5+d04Nm8UI/lDS8GHO
5GGv9014SqeVL7mys7G6q3goOEGFLhM4jXx6AwnjEuh7zYVNtnxpkFTF4fYc+4cv
6rtBXoR3qGA9rIbuWHXBcdjprW5Mmn8+bEhbnTv3OeHEKNIJZZ1JLQIXdYtfP66k
Tl5SLlsnyQHUKg6cBKcX0ko64tzcaKzBF2pBaRV1fah9q7B4HlAO9rudrlrYei5A
DabrZuH5K0PnRskea32XUaGxH5GIaX+RWdyeulxI3PZqfY821KI7+5FjdvAQBvoL
cstiqLFPeeEitYcZvr7RRGFeLyLOwu4VCkx1esgAKrVO6wAzDLYGRsePfzcwhMCK
FULvHlfOJ+pjAbfuKQQmU1UGfQpR+pVkAWkvGogEhE+FvHgKJcu2vr/tfReKgSZp
NReIS9CPBGgwbPN/lfqKXS7pwf+UoMUwyTIbZWVirEp2+6vFYw7HfvbYaCU1vF7R
WSeEjGlhuDvI0jzLmlGTWEunryDltVKlxRPOtKX6a/GunoTKMDol9V3a0xVOxEAN
067r6g2+uWRCnINl+TlAVdUIg66QsJ4qeuWnYLydRCPf/O2K6VjtQQHI6I8o4ieV
yNoFyhxGhh5cVvBe39i0aNG/K1Oe/LcZz81BaSAe1NrUDLXDIPT9WhQeXw6lAmEp
3aupiOezkPNCgmS+o4UgRgwDFWkjrTdO1TWNPvCeqj5BxzCxnYZfiOjBfIvFaGjj
jR2gmj4pj8jdmnGLiIc98TilvcC1Kjj96jwU6gPSOQkJnbCbhr2a/ISkTxeAaWgc
HjrPcn9rRDaAyMAln2CH+7w7Mr5hRITa91v193A1gdn4+86JRzuezE8su+Up5vW9
cdkFbeZUVn6nELW56Y+tsqHOIY9Ao98i/w22wBvWnjZUy0k+KEdmBzWtca9m+zHX
hBi76W8HIYipsi5CAnjNo6ueFDIg6+1qCbKb8CZyV91n6umjVEAmIvC7TV6Stnbm
NTE4eePQdI2EPBqHRuvSigZ2jaB9Qi7z2afd3dNFx8NWY/1yJIzAlWUhOI2zJukm
ff4KHFQhgYNNX4rXOERBMCSFGDckOhpHbj6Cn/1LbtODlsKc6uL80LILPNwnWvoi
VRwatCoOoRPUmYaPlxMQzjn+Kp/IqHGmwsjcNy1/3pKhWQL28oqczonksrPSRyFE
mzBLUYmIpF+qR8I5IQHKN6/Gn5nRgNeI/RlQ7zgUpyedMxSjAGJdboc5BzCfM9oJ
NKtWKuWAvNxEtPBmHBnr5K2y30aFUfLa+e3ePWZzdD2y+vt/u9DwQYNuKK82eZh/
df/PWHyv+rKjDexgNP/238UcMTLRfvKtVGqZR6D5WK5e/KT751VJdsOJePCtL3wZ
T4LNdc/ikLdm0kgqayRA69ulZVy8jWuJwId2ZfHXO8rw+vNBIuPcPLC5H23JUC10
j4FzDf1vhxe+hZh9Te4dcnQ+Lc+mqM/r9YixjywXURu9YRO0v/8RQZohR9tQHP2n
DfqpErMSwAaJqoX//6QNi8nR1wno8rdNDnODXRjbuY2B5TjTKji4zDL4E3ZfowzO
DphEK+0QQ/TC5uciFdudvzfOUYp7mHdyWs3WjPk8Z13I8K7Iitx3t3Nsg/3Is8K4
oAPlCIXp/rpXPfIy/JjeHbBatv+jhJfACh2laJ5s04T8m1xHyCOtvyukW1Un6RJ+
v02Obtd/1seHAu0McxcDYRAMEfecpM3FFsWYWMZHAl3VsgLt4oqkoVwlFQc0RFuv
tQ+v093eRHP2uIxtgPCdZcU+BbWXwjy1laqHX0gPfIjRl30CHgFqA1yTwF3J4dMA
RdrgKAHdHrK0WilckhHFRs5sOzaw6UT7uKdP2K9kxDC9PudMCQ63zXIobo7KbxEP
6XwYe0sMA1ACD2IjxAyPs0wQQCfFf9NJYPjo2IHRYUW/8yOXBvAFJO/24qzUT9RG
hGZOshLXTWEKGf8OPRQRKQqQuWwB2nd1AbbOrOrJEocHrniNXjCmCuH+qGx2G44D
lpEQLr2xLXknIAackQ1JHGibhYVPxABIDOEqx6jffHtvtcB8F2xZDR/xhpqg1QGH
DdzmKW57LeIcw4ZVjOjTlOz/h1OFQfDoHM4KkOpuad422dCy8ZvoV3AK0pdCmVV0
uiquGEIktEROIapzqYHaVUQpyjEl9Jdt4HMUUkykFVYnHt5SJroJr7eaeOjyXGlm
aqLnXmpZXvK5WUcK2nAk/cW64edFJXG66zU9qG97kCoQ7yIWn+peO7rXGvILcaZq
byma0p53+qVQWpHGp+4QHz4eggZQTW0v75iPWmIr5eFJAMvczlW5ynCE7vyJtdby
6NAzVjC15MtOYzw9+lZuEjF3SQD5affWfle5U3EnQbxyfj3S12JBJkHrDGair+ZH
S2K6mYMpPhANXQ8Fy5tsfxVn2IS0Ve9D/ZygIn8epW8FwqU+sgdY7qCGBsf8KccX
vFUw1QQ8D0Hfm8mT9RbEHXESujBs0soKul1u6GYBnLIXLgjKA5/SJVSF43dooODb
4QyxVVgNqfuULRn5hIZ+Twyaq2vVrRTUGe1/wxWQ815BxxhN5wDFtqlCo/a8pGLb
ALd8hI/8gnLZMaWARpKujDVRJCPXT7TffdQyCgeMYJPOkEnB116vGIY5tBihk0pO
UCkD3TntJTR+zErUNO5Bdmc/JJbky1u6vgob4co5SEWhFoE9T6YdsmPJGcOFJC9P
N6Pu7HonqueJvelHCheXa5VMvzHPIwCz8f0SiGGin/ELsWfKHL/looVzzM2ZGhe6
q8Im12DTCKILWUOJVnaepYsHPh2Nsd2WZ4KRkdhS52Lcl05ZHsG8VyyQxsT66NRf
A8rP4XYCaZ2iS9rcgF7cW4+QCydckzJ+mzg9TcbgceHB3Cv5VqjDDRDN8ll0i2EF
4DcZfcJl1LgRGhKmm+IMb+0c0t+kTz3hbfq4rQavppENxFSvWOhgBIxBgsEDM+gp
fwYb/Btf7qjncIQtuqdmAw54yKFAFQyfmJetl0hlTwK8FAuqBKAPB9wPMV/Aix6Q
cpnM/FeL5uK8SRBQ+6cUGmjwRivo22befp8pqb8bTnZtX922O/vqqcxAYx1nBQjq
riKUrMZ+FswYQTslICa3mat4N6AoQt0L3O0uICnv2zIbTs035v8ed7ykVRTDIVyr
titVvumx41tveapcKSA7MKYmnRlb1crfqtPlbgS2/vezsJ3sZ3zVjbEFrJE6EDwt
VBIf2vFe8fJfhv04pdZUQs9KBVW1qq6pezf12+j8WYzp/Blbc1/8sOK9/yyinjMd
urAdjtjxMcBE7nQ3MbwAND6QJgtx5kuZkX5iAYyscbXu7sIuruxsOcdNA0vwDgzH
Upp/+r4tvhI3a4bhGhLJr/SlrNb8r6rBAlg9PlS/CLroyx1f7kk3id5GqFbakI3R
qHsC/3ki4ZCyviPRiOhPSndhbbWuMNIdgZGVDNzhF0GU/jvEoFCRbOajqf1fLkMo
XYUkieLOn/X5pqRvNvPfCQJUQdBsXudttd7eSQhlMVHjV30srSnrnfSt6GdG+E+v
mjHe29tuJicChIA1c28dTwrjQVYtD9P3bkPUx0qBcUti74Ttn+pxpjJAy8NXYVFI
Ol7EVvDTtxFHnPnJ5zrsS17MpVfnkVUFUxg+4i5p5DlXzaPe9YXhYFaGqHDzW290
z24WucALTKc78FJ+VLCS412AZxwj575ndcNxhF3Uyv/RXwZ7tef2ylSeZ8Kklwd3
BbuhTiwREmcuyOwSONcjpq/j2oW0FHnhWQbD/xwV4JD6puf+q+4CZiQwrZEIRh2Q
JZO/o1NdxgGL1S6T3S6ykCy7L5H3pJMhF+xqpC/a6Ez01MlDeUmnMD3br72DeBbD
AMokUX9RsjriVEBR6gUinmjOBOBFo6emytjpjrR+FbcS6w6SWiQ8Fjyl0/YqamLv
+sYJ/Be+34lz5i/PwmsHj+XwnaiUhD/GivxYYn+v4BFIr7+T8RYMnhMqcP/TgbCA
5PTmlLInoKI8u+YlkozQW/r8fzIhPQoAjZoGuulX3fXjFdU0gFjA4Rbtu2UVvIKE
EQ5+EbiNgu0rR5SDSF7pJ7jkggL17W7klRvc3hj6WxtLeu1iOE/snFubcu+psbN9
PhKsvWPzHZpztFYTlS5fN+qV8E8oUeTfErEDiyVHTuPzIHJU/IZv4z/b2e6uUq+i
/Zo5ViGoNRNEI9/GuUsRbmtKPcbHjCdVm52ZUi5YFdcOGh7Op6mtSgmWMluf9rTl
7O4xiQZnwGmXN1HnrIl2QADtS4Wktmttp/raS+rFNlkoqJDuoauwtHFNdOoetX/O
MrFLaFjOS+2nYyivnKPasy37yUDevdclsiDuGfCy51PDNvh8CV6Upi8aJGemcWYl
VeJIZdCkzYcAiKPonbVvApdAS63temZeUsHa3+qUGygwmiRd81fmrlGlCYwUopYt
bhFOHIglF7Anhgxj69fZ1NXIjqkz5UcW1a/U8tr+f5qYhEHDeBbeKtw707kmJ9P0
G00rYbcgL9LdODKXPYmECYfBfMsVyTrZWYFROo7tLfwNDkhdYrFetRtYo+W4BrVg
UH5lYcDkhs/syvOU5txns2ScxDdS+YrioblYIE72Q7qoUCUjAC540jj8/PTzKFoJ
JTYJNlsCSmLUrmVjurhXmNQHl98Euy3EqgcTPvRuHMjA57JntM6fAYoSiNtlEWHg
bznpOCCxDBTc84YH3tr0fW4QXKfhFYCirfFRY51yNyFCagSjRd/8x7sHGl6IfcMH
z6O+we6hiMDM6mCggNrgPYRre14vtCshj+NE0rz5lZnq2pAYheLiBhwkjvRfPCOo
sUr+1JhYRPlawSOTIfB84LmX3v5mU1tv89+i7iueLQ2PgKltTOsEeJogsVKziJ4v
w7Vj4/RKGWWjJjnDsO74qU0VRqwsLaKdoMUQI2KAyJnd+c8/YFe/Xvuh2d03hu5d
8xtJ3Zxf8PTZTSLZzMSWl5JUII8nblI9jbzHWzCk88qkaC1lqwkqjiAnmNUsF5GI
mxIObaeiFBxIwR8zQG+gRdketH22U2jpc8WdfBVwYLcNE+byXUli8C3/L2uAt13N
UxnzXA5XUDzm1m3LO/11bQiSPiac6JzGPqmRkF1jtln97nVYLK8jiFUw+Q9u6bdt
9H8SFFxi5E5S6fF31eR1/YnpEkqAQ5MhdU7HGY/I20YjY03y0yeoNgqPSb499Bqg
MDWe1hANpxvenod+cpPO6jTa5lvFEuP8hyOOMkp5lhAY0rZmaU7/Djjr2XwbCNk1
nOvJz+DJilgWUJGWNmONOMyXYTLg1wvQiGreYTN8+k1u/ITTS2xntGnc1dVrLbxp
oqbGxBnXHz3HQ8iy7Yap+HQCBvRTXi63zvKSiAWoV35ZsJW2CeYfWbFyouuNF8s+
6TPVrBPL0sLKTxPJxoyB5/F6IYazVXtZLNBJIgDYnrbSWBYiPiDwK6vCwUxNLt6W
hMTm4qqlUfMUNkdbBMigVmK9S6FmgCXIwx+/V/uWyYf9RmNI5IRRI58NmAh5ljju
sI4OTE37SviN2OAGZMEeKGyha/uhuM3B3+UKgP8LQKPiFJdNe13Tx5P9KermCq/R
12iYX+R5vVXBgZwJHrLoDyC2KT5gaLtgfwY2+IJvJFa+GKMx1H/RZGjUSjtIpeWF
VdVS/RzqxTF5e5YYiPrrda5lli97N/IxaFgZ003qlcHs5rQNOt7/oF6l8VVsXXP5
sWTzu8vVziuBR/cK8GCIWORLD0rQq/tNHYE0B5RVhPXdKk6nOmaXDMwmihMGfYFA
goMl6lylmaZmKOzMmy6QI5bJ+zh/Zj4Wk9l8Iha2RWW/vyjTauGp//8fn7SpCwFI
x/H6w2VcNBeQnO0/8J1vqgTNKTqXqbcKAoUA9GLga90Xx7FX/H9RJp1C6j+TLBHU
e0YiYvnaqzS+iE3pRlUddbcov7Mp3nEKosgHevniEOsM4V/wfTknaSIMoN3bEhsB
H4q53PeOKThEiZ49P/27inAQBa8G/dlUML5Ao3WjyHipdLy0s+i7tkDlVtggO/J7
FqO0FRtn0z0TK435ayfTUBRuQfg1jUM+7fMbmNb8jAjxHjZ0eb8rGewxnbFFPbu4
PajlFEPvRPQZF8+aDxImmwmEGpZYgpJkAeCK0x51VoTAMFYmHmad67Bat++qdPa5
U2FsuSJX9o4g3r9A05+5oNh2kSnCazxt10M73WwGbYsQ3SQB+yWjZiXet6HMbE9s
QubJPQ3GMsVCkk5MVWNfMFUwVa7/xx93kopzXyTGOIJTNkHK2g62eyNnRtzTTXkf
fMLzEvZv/Qh5Vk6cEH38v7TVtkpAcMGINrIaCZzjkV7UvBcS2LFaDSjeTi1jjM45
rT/frlHPGKdw4GD+JSYHbkrGaIsRQzfKPoPfBArapuBVXjHFbBvt9f57EiyouLky
Y8aHLdrij7aGXcL2TKa/92hvJ7XaV1/rCSjGlhDZjw5rRs38QtSpp+yK4oraS7F1
XCRvU9JtA0Q3W0WQ7DDHtxV/r0fqq3flitFSnUGbWGVE8mCQOid671tNn3QswaJN
QvqPD+fzlWdmdJrn1v2+dvU3NbN1faldYuxP8SBWeqYmPXqav1ZljDofTXRj5Pm6
OsjzGYdxT45p92a2DpQtlpQ94CLcgDnEpcsCXV58gb0t85ORmG67ErzL21WdFfkL
cTt7IyryFOwhiM/z+7Jr7BhMCkZFBO6JOGK3tnEl58H/lpm5wAfknVYJByc3Iy1b
FS5NbsBU8nG99fMbeitWpEhOXpKo0bjjitsp9QhTwYfpMi0AvuAL7oQO/0Oojdi3
0qzvreS4uroWiXbEy8PsJ7fAE0bEk8G/WwLXmUKbn8faeXHuqNEIQac8uehEcwgD
L4eAsZ5lP0Z3HK+tfiNUci85LIQEt5nwdZbpAiOleEbeP6dM9ZfOMpIwy7b+duLH
M/LOtMVcGVToTJxelKNsMzvYAhCGZVcgiPfdOz8MR5dV5pphf0SRjW6kvm1U9eEG
aoIPOkaD3Xbj3odcAxct3hjVpQRYk0/vlPMzhQ80peVZ35O3338H9yfot/ZJ06Ps
KMLsslfH0vig31wYPDUUCZrgyQAd/+B2W3O5YM0uY5XYWwpFaiuIVM3Jk2DytzqS
DRojvELtq/sxK2SZfkYXS3Yi4RjJGNTThabV35hcHiJjWc9Uwvo15ZjZpnsyNMwq
qQrc7XYofol8J0rFmDO9Iqhf9MPfHeskhjAGf0NgX5EnvNGUuKcsqk3u5SUJWgyf
sDC/gNZ12DpTmJiE+uiZxhf5xEJoBVZn+c0b6KubOCaOI1NnuOC8qCzhHlFSOM8s
gRZzz2pwz2qxXtLSwlRQRuS1eltl3X/6YebyoMh5BMLNtgGOmPATVg0YL/6gcBMb
8fdDnvWjc2etyzSA2vgbNwjzvaJgb/HoKw6JKbht4Z4zhYafpDa0z0cMPoJQUbfa
HvK8aBNauj9nvGFcW5bGbr+qLeYgLbrgbrQEVfWFoWIhqkQq67xO79fzjy1XkZsG
WI9WP7Bo7Pg3EduSL5aM+ZvakZcNLmAriKy8hkQlt6N0al7o4EqT/o55R0KtQJjr
jRRnS0F4/0U3ANuJ0ux+t9QnD0BJn/qpmWp+XVSJM1AYcLxV8thslHQXuaRmB9+Y
OFj/D8dTy1nzPxj7WgEjX35lfeWFfRaBiLUn7I9v319XCMJESSwEfewOCh4/0eZ/
dJcWX/RAzAoThFY4YHiihb1oe1wgL99GZhx45xL9J5wXbYGDLfwTxjsdpum/QU5A
L8gpzuycLC0eG0mnfpoJxI0yW3iUxI1PNQxiAMw6Bw+M79fF/pRyYdYL2Z8rZhq9
o/U4jiA/gVATG2nhG4T1mazQLlQxbydCuG6OZ0csOOI8oKytZKnsGmZ85HbaMWqs
+wwJbaDhFjUERgsWuzkfNGpmvpg6K+xCSSaMuH3MmTKufyCCqLY1vucF70LkdBto
W9t0G9yLVTflm3+hMQ1VsmAukr/J1m4/tuMkHLQmwE6eJs1usktGp16P+1Kko1D+
W+HJwcV0/oDhoFMPpKx17xvnu8FQaDPL5cAKuMWHUxzImXJeRj7UtDrCvx9NL7FF
l4tnYi+xOSlPwmZOlswxsKV0CJaCBZcEpwR8TjlTRLARZz1VzOFClAMi/ca+0iRl
rMZ3429PJPEETWMo8+ASpcAWXMj3diXmQTlAXkc9I4rz0o4ecOlFm+barhK82ugj
bQ9ap9bPcadwC8TLPWs1DObPtfRqaVNAqtna0bfxUorGO8tYSxuNf44ovqzJDLNm
cNXO5DKcXheMLaJCeDDH/i8YOXZKWPC5hCWm+oy0KO9AxRKdPnOa6TYnncsCVkFk
GMmOg3XaHzaN7BoU47uIlXGTJqTNwRT0b13+M1gTwV/tg2hY4XurmIJJRNzbwd4h
+UUeWK9kmCmLNeEK3HiJ+6TmM1nwzGuXV4ZG+Oke9WrlCB3bpFbpIlIZa2S7k6D5
kD2vEBLaVunDwz2uDsnZBBYoM+f3VSLwVdf588p5oFpdypXQ99phblHE5Kr/vFL4
nUY+QiHCrKU2bgRdVGzPP4SC/8PgVnrgf5nrUOQJntbEs6qT21SrIy1sHQ9TyamT
Eez3+dufZgDpVwRpUB9QgkbWNsYXnsji1rsQPXtB48TClflhRm+WFjG8kQ5F41sd
Wxwrn/ILjv6vAMwKIvTj/0cf53y8id8EzbNzOIP/540z/Thdh8VOQG1swMLbEJHH
hRnszy1fsT80a884D9+II/XqeQ38QYqg/6AkAV5BCbT6DIzJnoJPTLhSgT8DO68t
RpgHBTUqr9q6B+zON1zx+0M6BJEYMUYCnTIQzSaB05lPRLZN6TRNAvYrkd5CP6mY
5BwxC6abCKlPw8tE5jBWjzRDoEDV0qU0dsk6PPTGqmfib8qFhTfHEACD/POx2+mi
yqEw4HpSsWng3TtJDuik9lTA0XcJdgDHmmqXLdlGPvId2z6bJhj4zZ5FOLSRhKi5
s5MetEIm7kCIBJd33+R5QtYgg+Y9mRXl8rp9vMPvBaSDjS7tdwZb0RTLblqsDxOA
FwZc3ZpGWhvXiqwtByZCD7Z82yV4n+WKR72KZEXWXhGR7LCz7ybdiLEV3WrEnUzV
F0sARlhdLrZLG6J1I7310nCMtJZGhc+JOe3vkg7Hyaw81NmR50EzjDbZMhN77eOZ
q3TOaXS4oAY7y9NjvAqzkpum7JfI154JjabmYLA2U68Wswxwjl5y1rREW1Bvs0En
CJfil65giLINLp6VJyraC/nzOazAATh5bYauC9nFDItcJffJ7RiC6BlUSYZ+aFR0
oR0N+jOxDxcx0KA3wia4j6Kjgdj2goojsnB8Y4K077b+J8hCBUpYq9rGEdW5azkn
q4WJtuaAUHRHYFwIjJZg7TGvEkwW86Blpff2MgMc0dDjXRduszLFVX6xL9w03SH2
cc16DXuhOvUTCzrSUuXGtkCee5U4F/+P6IVqPQbNpGljyVVHniZeAA/OjXFItgDe
iWAn2R5IrPHDpmG1xIKXZa30pTcjcN5s0eeZgWmkZqCgsNVSedGHMlrzQhgss5lO
t/XaGeWefIJN1wm+KaQDpNQfE3kE8f3pL6u+nsIglMXw23YmzT4DhxP2AzUBtxGQ
3Ybq5JZZbcfz23zIaGT5PFAS1IgFcrVWL0sSozZ250HeJvwV2Uu+hLw4m/HIwzoh
WVH0httH97CHgH928vgEn53ThAQx17dMY3ePyzJFbPUKa+jY6m+pJKCAdbTjnZUB
3z6Ra0HkoqgTjNVpvRe8XU755G5aGYOLNZcdOeGmhKsQtn4fZ+g6mE+SkLFJz+xi
67oASI/xlnaUr48r7QpucRyJJQylaGun23K9UdUS+i2cZD3aIbOwD2rUrUaPGfGN
MEaFk22dmEWKkN3v99Rh/6hmB8xX8zsiwFUIiPlEBSgQYeakbLEb4fz0BsO9PAxN
2UShNPKBHzWAVt6fVCh391bmIZLJyM73CpZ+4ntQmT32NfQ9gc3lxASLyYEQ9Bx9
9gyvav+HelwvGOLEQFHUwOua1MHyr4r6ML1MC/vFfsizU01nxs/BhcjdQppSsCPR
lAg2GrL7wazyK7l4gD9oIsrMahrP1TMRgeKMcljmiZxle8ji8WPFS3Z62QHT5MpV
3UARhUC09nQTNjufq8c+/T8h+FWR9zKfrKoN5LmLjCiZWGsyk1y7M7bTCBsXbpZU
CQz2ZfLx8bEqBmdcQMcf3tUSmHP4NMX6Lzr1SPMOJ4y5ji2R5OHHBswawsc7tkC5
+nLer+HoBL0g2tTiN+4Oq5ksmHh/RNpkBHI1cx4mXCueg33E4S2+m2TvXhRmoE38
R2Ti05PbU8e2rfx4sZKAPQKmZiBTAlsyhv+H6tQuKT8z7gjG/TqpqkLHaUFmSlV0
sHF1x/RFMQv48Bg/qtSiiZPrKpLUF8MRO8gy+JZy+Crn517n/+LpDm69raIRCiVZ
9nzBQ1KcHTh9/kl63J6G/HYnW6WX/ArbGgoCgaDjWkMCVzes1REiXnvLhBs0Al3x
VJ3FntirUgDo+kh2MTp6jKwhV1XvfZ9X9qBFAiL1++hmDIf5LiNxO0c+/j6BOazx
jSke+M94H9I3n8krih9Ds5mYMDnQh4ujS/b4CF2ivkSxvJlN/SQKEdtz+yUVnDoS
phv138VOfB4N2QR2hDIA91+1XiTzUYNjcfA5q7NVREsamyNXfIGb2h+tDdal8bUQ
4d3CfUWB213SKOXEcqP1McUalw3V7o23Ky2bpp4cIGpYBJ4kJqFE8XN4STkP1U0A
DSljOyUgayrbhV+qLVlzr3lu0DIX/YHl/pOwx01nI5d4zWe7JqymMv2FfB8zLo3n
8fdaFAeVzJtGt7nYByKwzcxKPmVJ39eUpFSxgiqX8ml6o0gMkc1zQx8HuAuCS7wm
r1LyS9I6uzI2o9zOZDfAazkkLQBQzSKMoNctf8wYkPXW8YLKzR0pdw9F7+OfQPXS
d91ZL4FyADQHjUsO/HtlCM3epRmPmFNequ9X8AT5KxX6G8SFff8T3P6FgSTxHqO8
ecss+aPaWiudqG15EdY/vvFfKPVJtHVhE92lZMonw9n7JPJxjnP1sCp6GY4r7BZU
sDvtV81zbB3QEfn1gCgSp3JPcG2oqr1GMBVNnyoNHnUbFZ2qOcklbYqFGcr44Ma2
fRz2pjm8CzDiMNFj3rHEIjgKnlDloupaNGgRi8f1hDuguNr0+Eox+dlf4O2WT4rk
yLPfmuAYpm8Z4eHUL3Cj6Bf5qt/ziYCI9hh3iHOyd2TdIPuprirML+tykrQTHLsV
8gO167Rnxl1FumWy/JLbhXOAO58pbQZV2mw9B/3SwZtGaFpIAdK027U6uEs4sZi5
6MFCcblJ5kIPiSV5snKO4YUxpkDppFfYURQYolvjmWC2y0mY1ug/jeyfLIFaVS43
NAi+4FIDQmddQbjFUwpOrwQz49upL3gWZvj3GPrBtFlOz2nRi8MRFo2cOFVIgW+9
hD9aJ1DM8HDKaiKI5h+Lt2kqzVK45VnHhOiG7q8JhP+Jf143z/ktMU/d3GM4e1bg
GTvgyNtOumkeWE9VL3+dakLPhRFxNcAAUJyE76aP97TL/H0pv2wf9z1hBNc5xN2P
g13KL4wK3edyOKDlz2bcavIeLVIqUY1A9B4+ETKt6s6L0hHSEHPdxhBiZlrn7t1a
ux6Mj6L+cTYks8cuFfVkpr5JbgU0y+UcsgGqlbaKZwqXFVqGrEyvTZ5YFe2VmfZR
YRFvp2dcDYULj66IIDKVSeIAtU4wBDHcSR2+iIXCHGPSL3PovI7hhdGraeR/63Bf
vIwqdqIYZWuT0gbXljZ1x8nMc3Lu/W7OlpZTsIdKNb7MwNiIWTCObwm1yNRe3Il5
i9qnH9xtiSsfR2G77UsUpIGdJJLW7Nr7TkWmfqZe5R+rS/pLcNmzGILNQW6lag70
DnzTIw0NenCpeGtLs+4whcsRkJBkIWLFa1NKsPyCgJN7ykQooS9v221LDzn2F8e5
xd5dtlNmJxNuI3RL/387eu+1XU1foYciplYWaTXobfc/r1yw+BQnGQHWfhOZFiM6
DRf8G3iSBOA0uVx9V2FcwIVPyyC3M16OZdCKtNplnvIv6idcaRD2gs1WDaKn01bj
zpt79H5JCGGO2NAwTWFpfOBaU3uJGE+Os4f0l7XHSP3ofIf9V6P/sjf4QfT28D9x
VJTEZTqgeBFzM23b3wHv43FufUIdEfbYNPSKAflU2ryX9F6ZAqtnAMwiUuedtL43
oc+2QFm/DPLli+h7bra6civRiheLI/kLjeCUoqbapVUKVrt/REKeZAl2kYL5pSi0
z5dcWBGDg/XDrKBrLGrbm0RCdDnZZuj0hBlf47RA+uTfdzWWpQJ8GS287pMeaeVA
/fbl86ur9QKY6lcMTnhVscgrWY+O4gn74PIB5GBfkf9yXL6LnANJai1QQjPEWIWp
YKoUwmdwwpRZvpOmPFGMw1yddB6X4HEG5058a4ZI7PJFIzk1o0+aqJvvnorxb7GD
8Ehp7EdWDBWjcyWdlXrh/6D9I5Snues421hukeDYZ6O6PssmOeLdv/2eHwHW8Yc4
1mzD9R4Qjy7NKtDk48DUKBwBois9XC+8vnoiF8AuAQt9cPoG22JWacI4tz2JpyL6
lUUqBtCZv5oiuPYGkzfnxVqFKznEqpmWnk0r/GdFbtTQnvcuKx5g5WEDDqKR94Kv
CVErgOmmhvvKMqJN6WPMm4gx6uUvFd+dXtDFyO1tTe5BAAy46/qPperCosBXdFLO
XrS0vuNBNhXSP/6MBYPZnEy2OgWJHfLHR0MzXR/2nnLkSpCcvJRz0W++41hWWzOe
5s9iojGQ/CX0M2qaXTpJ27rIFT6PFAhOvX1y091RbteeWUhGInPlTRu+yCIvC5/N
QiCIC7ydTZzijHyvcw4IYp1h5PazkulLp3F/0K3cVCHW8nl9xj79I0q2Jnz3oe7v
l42Bmfu9jCuM0YY1OrDqvP2DlxtQnnXtrgMLQGwQW80F07rjDEhJBH+26dUzRNFE
MlCrsZLOZJn11oO93ieXCN3rUL3k/hg9XF5PYJcUia1eDuwBH6+3rj8yTmQAv3WH
QCKHH4NwSrv2laf0xmrLMuoozsbOfMc13WI8kN/nRkadyR0DHv3anaVAFCsccBwu
H03h9cHavhiYoY3vvv7KCCkSzbFwf1gqzIxfmHjHHOcuHuBji/uvth27aro8ybhH
OIsq0R7KAO5j5znw8HRob2oLtmrvjVGDe2YDmBCJXgriU8mfHFHfVtf0W2D0qiUO
a2gDFHp280oL9mWJbQvEcq7gGGP2Ms9GJ35mC2BNCs4D3aZxCYfNl12csMXg4+P+
Nh9n3iebOnQCqZH0QequsLfRpbWqDOKDUMwbkUva0eSJ2ZzNvxFjMaj6XS4RMx++
M52CbrTOThEM9dHmv1Gv938JkagIqBZ0OXkProcU7Ct9Th6QxQltWQt3H7D4lHCX
rUL/kKbwJc1UU+zmOmLf3oeaQMqWNyNMmIGrxfyDY0G1pRmnMU4PcubKUm+j/32b
9+J/LgYpcsktwO/cANb3cjx95D0whaQQxdxri660QG1FllHBIK+bojQJgRojSn4D
vq5HvHjtt/4e/EqOHabMeouzYie0Yv0IrTmE93Na/MLbN897Afjz95txDGRxVcwu
9jFbv1N9Z6ItwuqEyDyn1k9ogndVEoTv0Dkvf/k9Fw0bXdBmAzqCAqeeqZA32GJd
bGUoVwhul7FsELX1IgyOWVlfAltMJDYM0fMJa3iS8pNWoZIvMoLi5yrIdFFEaLJI
HwLHhoK8R0M4E7tlswK1ECOt2kQwX6iXKXfX3PHuDZ0Va57XQSS5ZbTU93kQUxQq
/kJCuEepz17TIWgoyVe1emF92LVej2ZE0thaBVoquVFe1gjp9FzRBq0EfMwRYrWW
yVOjXcluNvkf1PHkSIOXiQgM1jIjM32gLeMwYz6YbtS9Lo+qoMEtQGgXyekdszMf
lxyKBopJUaMptUIxi7+U+r+WZltzVK8NWfKnKDicJVyMXAennwLvQLe2uHGXE6YJ
c5rciyQQXgIVeakhsDAva3HgydNUU3p0/r3gLSZeSkHsLDPB9mnXGyyuZbE5rbvw
j5DW8W0aabSYkVSDgdOEZlK+Mm7gT/0mcOYGWtHxKtkqNM2S2P29ojVdsUVvDips
mfude4IIJpfa9CtwXDhHtczcgBj94dxKGlVlGz1Q7vxdDsyZsARUOKOowH7tTQc3
MQwHUKQsyOD/D9QVcqEZWKCZehUiOUiYFq1X2iz+vvVEaNovq/bOe/wXJGkt69Fi
FpK0fXBcAOEo4ATKdAEkcSl/vzSKYpOsa+6A1LSs3R6a4B9mDGAvAqRoF6O22BAs
KfriBjezEPG3Jqv2BQXXswhSb9vXqnIibkr8c7WzCSWOKbkUowmwFrv9GfDufU+e
ZZdLLMH91zdR7Lw/vPoLYlkcMXKv2ABUBnGMB9aoBIG/MQixEXCnMpncqzCPt0Ze
q03ymINIMD6zP+YMNLNU/yXq/qvk2QahSWrMcV/qDlf7ZmWuRSUkp10EpXYSPBiy
9TLqVvPCu+JJHgcaQAWmWXu/+INtamkgqtm1C6nJA9ovWYmkvM8IunYYJeNZtxcY
w+lOAG0Fpy01C41kDeOdkuAQR3N+4eRP6Cp0dc7p5JZvPcAbRkoOLxbxoIVr3Xiu
vPxd1S4Ufi9/KRyeFkHAORNHg+RQgRiJrEZcBZ/4nw+fkVzZvT8hRE370m/f+IdR
BbXT1U9/mLeM1QNV1voANrPKzzOlvs3XGYKUTYazwOF/onK/ozZjJN8btIUp4E96
BOz4qzG20geh3g1oufa3d8U3oFmjLkQkrvGkJo7b02e3TygIcPAZROdJCAzksQJa
GI7GCLkR0MlpwxWVHS5aToAY+w16GaPbT+JywC6RfhQv9/xFW/IP11ANmB6Xy0t9
2MbFKBwcnAffgu531emldJFY8GY+nEi0lAZBvcuWHW5O/jYZKQiz7AbkNxpyu5SZ
AFhEVhF9ptm5xLopeR9narg564xvo0yGd/lMgjqtV76rEPLLgBmumNpeilWRYxnT
H5iqMWMblNV7wS7m3RYWOZPMwA/K000SUouuVkVa2fsbh6dZsFXmd4wK7SfIdjlT
TESrf/IxJugTCzdOL9roz7SCbS6h9qbkB4hemX/rjEWdYIB0XFY0XBwKY6MV9GdN
kPJaCYfEjcJXLYxyrht6kh8BPKa+puVdcHKJmg0TaXjQxf94agqsHEyAoyLNgz68
idHOV8JBu9HRDFVtWQNvxNudwiLeRhmsekJGI8+vxmxd/iJF3/hV8B/tmqtFlHa1
JH5M/vGT3XwRIPBedZFDp4eYBk3oLL8zO7aIN+KPv951eiO0GGupNGg+ZdKyUv/P
gIVev76+AcmuecYfbHChcRnoWoLVleOyrBafzZkHvyKHnuvYfmiO3hnDDVzHl2aH
EulvGAkcJy5AEjYZm1kBH7VCQFNGrZIzN1EgvgQcTst74Irs6kyUKJPWtssYSffJ
XIwCzzkpYqXH970+yKUwtPB2iTB00ppSQ9YpPNfzlwvMeMxv4Kv9sUizMGnR5PA3
NvqHKu/7kaCdPg3y1Lyc6AWQQTfMeS5jYapt7y7DunmQz7MXS28tbMy9ysz/Iwi9
xvX1Jq9BuxLUrdwsN+EhEv0wUKp1rNqfB3lUXnnMol4s6krTycSDqkUa2v4Irk3M
3YkGdOMdpaQWlLbf6SMC8oxD+jpz8urTIEu795ynD9AjGQG2FwRrG7Lai8bHImui
bSEvMk6RuPtQ7EEK6EahCqgD1nXEtn/Y/QMDtozcM+vMZ1dGbMUgq++rZvCzs1xy
Ik+SBt4DKnMxkauJXJiA8i+VtELY42T9+7yP7kiWApo1jLHX845mPmbmo0pDo12G
72f5CLQlDRLgIDxXnZWTDLmmyZD6xPjemgm1n6Nmc7TXhg2CtuDzaC8urrpub0SS
UfUFkpXSN2oqygM8rZ422kfYjRrcLMldy8cuoLKVAPmpOSMWSeiMIPOrE3NVbkVW
r208qPGr/8RRcEFlUc9S7BvZG7s2yHgudeaU/VGa+//fvPyZOpyyp4a9KiKODydY
CRMhhjaYFj3ZQOQmMmJR5GqctDVmgJpthe9nQ7dey9+m1oankmoqnmNQztUGEQlm
QkA7sMoywVahV9n8Fj4ARA6x8J2/8OjD1pbfe+0j5pk3YKE+DFjrOLT/3g96ZNql
QSFiPZhZUg/SX5Em4/rUjFPOyNM7FEb9mJ0BiyuibDUUxMPVevsPUfkDCIveABn+
wiL9Scw6WtY7MobpRi5U28FcjT/mwbyJPO1I1FmgIrw5fopFIUuJiTrR0cr6nUjb
aeadOGh4sK9rKRF8ZWvKBgRS7EsMZk4yxxcSRURIebHG2u1q5kayZBFWqOKSmEKj
pJPp/yqAJJFQ2nEHhJt9I/IrQRfC2akFxDhV/Ng3j0SC73nq7ZEu+iYT51GqIbJT
xC81KQ1yRCTPPbVjRRPKgXwDnuoZ/CNxliSGbvd14tLXkLQmjnrCIlVQ+Gh/WDCn
6AAPFojZVs/UN0Mk0slsKFBZy7pWNExRfAnKIiugnu/MhGlP/5NpSbv1euh6HU28
nF/UUSBFXySMzzF2bJ+zhpus1YaJHB4hw9dzphVSG9zo48H/CiAeXAbhrzHUUOEL
Fggyofb+05LJTy+61lXRYfU16MAzaBG9AcmzYqUiHOakhS9S+BS52HpuuyP2N15Z
MXgBD0J/tc44apdrmtUI8TliuHTEL1omTCV5a5qjc8Rgv/m21mzBNwz1nq0kzl1Y
cror57R94QKlbsFCd9giX7ne7ydY5CtbmVRhoztOC6enRQEwBwJAs0vpe++lw8NK
4lNQO2EHBxO75btHwQkM0NRmI2uyVzyAYqhnDIdfxhdAft90afRK230fIwL3HsfB
HD9SkjTcquIENVzgI/KjQ4sH9fs22jn3/S9slo4CfvwD25zUnRyXCKSYP8Eml+Rq
yQ84Se81yk7CdOPDCohsHzXVjiMB/R1PtzKl6nhCsmgXfCxLrSYeuFaLuRHRvlsa
rTYWI/vO4RBZ9MTAcsErk/AUwV1WtnCFiai0unohvbsyTzgqCksNk+77StnYqQcv
26zM6KT6RrddQjA1gMR5hs+B4U9MKdke29iEIFTyhCweD9upb5YQMxmkuxa5ty9W
qB84/ynC5O2b5E9yOnkx7+ZlzYarnBOxW88nFhn99E18Vo27Q82oyFDQ7+KeGkVX
snz5QfZim0FwvCJJpFtYvB+Dqoov7qpf8KpM9lBiPLFb4e/IXNIWGRC3KGZnUe+4
593zOD0NVa3G5oDnfTsdjtWeDehC50yiemKcugK867e0+vYhvr2YcinK5/ERIRjY
ntmmj4D/zSNRUklivPw+ueP2H/lO7qdMbY4vnp/JuaIboQB4jUNfZSXo+4mZDlcV
yRvAvsvh06OM4xoib1jLn2J0c3WxH0V87p31MF08HPgylUROtfMqrRNP9OfyJ1vI
1XhNpKapMXcBtpHKXE5sXItfy1eeu4Had5VnwkC9Q3XJlyw+6ZCavGuWx1QV+RPT
PPNphwseWQALjIzpKu23H2uAhHSfArlfvtNtitxsFLsLxqK9NQmg9knMKwx/tXn6
IFkKYZid1dRvdPfHMLRXemZ6fCHoYKxzMDawnQOHvcXrNjqGrbgYXAp5C5TO7ERv
IzMUwpuFQytbpn1DDWn6TfIxnJ8sUXea/MUE3Zt/xmBxn3QjiSe5bPHDkJwxnpdt
NMUTFEglI+4YcbBD9v/uMp3gXH20V5qb+anAsEofVg2YfdzlvU80Yk6I0r+nonR+
n3zOJRBvwO622z5TIW7YGLTl1JpnSvKzk63xXZywCJRIjjxAf4052mzpVx2IWiFS
KpI7iVCf5cF9e2B527/Kag1/Xu9ZTZ1+2S8dYUNRJ1GpUfPkWSZu9c/n9ChO/wjk
LgFl9fmM+7sDCuMChD/w5L9+ite8wn521xxcRiUw9Dg0t3DzRcUhwpmM/T1cWanT
7uzQ3pJK3qXkBcZv7QnbmNZSIWL2Q4ZZqmwlmvLF7kADGMLiC5jefAPt6VDeOQO7
NQnv22S9WqzxgCtDehBNDinND2C8Cyf/fJo6oicmNtNfzfiaqwQoiw3/vEj6Z6RE
DSa2HV2gr9VOSWCYCCc44QP8dUbihCUBTQXq6r+jQrCZFcekl7TbPp2/maV7RI3M
BCPXVcIYPDO7YAm2NHIvIC7/zMETzoQV4Gs1h//cuVM3k6obsBDfMgkzwqvRfQRb
U5YSyT32Ng5yOXRNmWKukq+zr4KkJ6AExLCVPGHABzNZiwPoTDXu+aaCjkQVMsDQ
WuyExgnBHU5nvIVQ19HqMlCyo3jW454E7FgwA6hHbrGp/zL4mbd3AwEjebTAO06F
O1cxVhroWXrQ+04ZqR/9vjbc9SCI1FUD8VIMt3L7zlXKzIf4k5X+Yrx+zuIMYYUL
iZ7towdlp2BYlXlZTpgwuMui19RpZoa+K/7Z0g1XgrQt1mcpKMKetg4PQzJfsztH
hD5mVVsJMviRvSNjQQ/4JfyCpTdGBgt1EOYyp8evy0rPuKwIgvQoz9a6ohacFJph
D/oXxBUoLVk7jxgs9SdzrU1QA4+TqeNBemDGp/JbaQ/8SwrsJ7dbFd8xx316LR9O
UG39hxbwUBAAJs1dOVFs8XGkuSoVQbbEVKqfC5bMazfN+JHsVNaso8Gh0FZwetUM
GDT0b+v84r6fl+P7D/dm8Uj3LUwhKqE302jIeuZJaeGFhiNkk2wbvmIjOhTnhLg4
SYG668UJ//CLhVUSgiZkBZSIcLj8lgKy8Oj3ktgPUYqznr1KQpDH3m2g6IRNaHO0
LAUTacFKw3rdPO6reatPLfdiVdoa0DD7YLQbqOeOsw3V0c+sQNiXeSXHcaayCefM
gklJsNmTC4fGh9EGW8mbAeSULVxt3cmXMwKo+YIfiHLJFxHEH2ClamEVP7P7jtnB
mMDR8XSUxa0IWY6bjMBcdJZFdFqi80YIwxjqmcDOCfuwkk9JKTq6VRG7pKnU54Y+
NsH+KllLJnHjkaFlmbQf+pLARqSq/IWXB5z9JihILjb9vy0WHmrBADBz4kdQU3aw
UkzFg+iUI4rIA5/yPyV9iYPTJqI7lU/fHjf/aJIWwPAQOIZ+KPHjPQ6oqRfzbgqd
mQIEbYtaB3hzVJ1ut0CsJRYR0d/LiEFZMwlNUKf3zMnMIJggjl/C+Yin+ePgE4Y+
/jZdEVPLCRTpUahPgRVoOucmcQglXWX2OOWBWYhM5EpJwKIwf7qqpRpaLo/EZ3qh
8rUNGE8Rr7FQzRM2/wRVm2GL7mge+vlHp7+CuKHWVpW8cwfKWgmVlBuhlEEiveGm
QkuUhRBkow4RA438bg2ox9sszQZIwoQso5xoY4ES/b9hjIIENpbvpSf9PYQ6JEBb
Kb388nnRLDFgAVBGGigBffdCF43+pD9qapi8KMx/L2WRaJ53XmtzrjsvtMPe1jDA
qgC3WS7OsIzMDaM/z5Y4MpuuDrqgpYzMQpafWhzPJO4ozA/48e+ETMXQ2VXQaxUT
STsc9BCK2d9adWju1jt3iLCH3NsOzeAoH2TXZTAASDSScob6fwqV6ZNji7twVaya
nS3zo7ll2ecQwHh2sMTXBDq4xi/MhGEycx9iv8qg4Ts+BUX2Cjedu5K4sJRX1vki
N80Tto8ObROvSB/DGQ8lFGbqC6iWcdDBw+KNMXEdGlSTNIKZuncXTqsQiErZQ2tQ
ZvLwXao9g6Yqp+VblTowz4M0MzI1egQ1d/Yk/4CAYteCV6frdJaWERbm3bzS6c0u
VXHE6GhSYwIlnA8zCRC9MRdTt6Tpx8/yN6f2Nmva7eRQJtStIMZTInB/jvIGGJXX
NKmS2E15PkymQNPFnv74mrcr1//bIEV5C1IG9y9t1Wt7XvQmwn5k0RSwALjU1/yx
EKoZ46q3dtcy/x6+z+DFEFvwDYAFCMXFoaeTeVWTunlCIU3DjGTgFcRzKM+XHuU5
NRtX4FCV2fcCi2ppMnEBWjv4CqIU98jEeumieasv/OLs5vcNKLbX2BwtweDF+e8Y
WGKBsPQgEjyaXiPUJMYCLmlFR1/nsw47wBPxhcEh/IdUn3UhAbMKaDNwd2RjWsD6
dOZO9azenFLYZPaK+TaFpw4p0dV7N8k6potaaQ3HUoLm989XXG5eszR8KKvhXjTp
p+VI5ZOn5M76EDqvc/BOWuQnzkraOI4jfecFVAXD4X8B0mtEQeNZiPfsHOb8AG+8
WG2S31ZkX2eFCvWrurHLEyfIuTaVGEiUMutnVY2yZJnDtqWXpz/4uMHmYFR0Pk/x
QKHtQi2ur1aeH5pTTfEmBlsHmuehq9Km7QWQUUIPn0xxQJLnaeWv25L/Zg3Gskc+
w6Qn6MacVTDbFRaX86qjwahJQtuRPZTldy5XTqVa/wOZFZbI7RtWFS512paVP7cL
tiok8N7cWsKNaIj5nUv0Y/p+Jt21M+Ub8Nn8+3K13TDdcXWIBxcO1UJtTyKQRuJR
FE9LsC5ewePgYSLglCELLKwpGJJg8K/HhpMd+cXZpzZkg1+ie8zTq8WW8kVO8p0n
gcxNMRmCRuXZsAA90dkUu/qJqdf7sdoBTKClTHwNFxTEkYErEL6vwu+C6/UBv9cg
JaG26om4C5UknOIPAWxZiqGGfX9leQ3e/2oqc7imjA67NaAxdtawu6BtxQKZ4qZC
D1mWgj3Xttjj60vZ5VlXNrJ9IsXdGgQHqy+YI7wZy0e3TOMJQwdg1EVTos8Tcncl
eztbewBA5/7ilmPOB/1rCSv5wfGBSB56otAYNOuxIeflxwU1xeuOqPb/i+JXx+BF
rIQLv6bk3KBtAJjwRhHzAxeLE5l8MbJMYGeughLwIxLDA/CF67p9gFvQf4HkZutt
OUNAMw7z96YY41BayPDviyP2nABh/mTqZb8DnpxoQBNxMNMGYd2ivBOxMXPexNVP
h37ABOvI70YL+KkusWoYQ83CK/bXxGkP80t+4AzMfaki6lDld6p7tscv2bdHAl+V
kMb8R0K5F6c4eNDr1zemml3jquY85MeannB1gTRSlkeSP7Y3q3gtfe6whn65CtrW
cgRV7HZr5FV3upbmUMG55EetDT7XG1ht6JgXLB8kWYoINFIGF29AWTQhvuWS1FY9
oAYpEerWac1JeejHsJRSfmDn5S33v+wJ6glSHxVRWYzxqiHV2X57STf8RyxdSUPX
nSgUsdaxS3W7cCK7//ZVIa7Lig64UjnIUnqUC2Wo0e54NmKm5cHr6iYMd4r064M1
cDkR20FHN8JDHwxMzVfbO+LRckNl9V23tuuQgSGd9C0a7bScBuBIGOZy/g8koi5G
9lTi+NXsZ6S4lYT2Gj3ogrZicyu0r0I7aLvbWOw//4cVmAH8VUZAninVB9YB4Ze5
ca7oAAGlJXQD1qf5ITROmeN2Bd5OpBFxSNUcf3mVC8MBPZvrn8hmiK9+7SZlyU5Z
8iLvRoSXGZUSx0pqI3qFr3dfjeGB9757TSD6i9CyC+1xwZhz1YS5vtrmghIkRc2Y
PjFML31gwuwPoxIJ/L97aEv5UyY3wmzTildIqqCGv2xHnzVWJtMpKD9ahqqnyH9V
TrlZEp+fqAVPjTTeEPLjmPt6Ev1ZU8KqYVA55aU/ck02cY+asGdISjkbhTYFngQH
ubgDO/nUpYn4JIipz052wxs5Iw+8FxJN5weAp0JNtL7n41IkhFgL1okEIJvq1Kcw
N4A9e1LyTjHvIp6BeHoe4UMm6bdCO7mUaP7EYErsx1XKwEAMEqCg0WMdSRg2Ekbh
Ul2eCRuoshW0q6Fxms2YS614+RDzWTqdfJcu5U7AEcpv5mGZlz8iMGQRoj5wkT5q
EV+8Fv0lezi3ieYKstvMRuBjUGAAABak2RU+RC8evF98Rimwtwc/fE4wymN4oxDB
yDze0W2XgyaHu6PkJFNoFz2Bz2l66ei+0rRamKUvgZMmpacbDRpF5N3jTKv14sws
a9Wh/txpdGcs39rv+4Q3uI6ZxwUf/RFChKcC4/0TD4p1oL3i+mNVftLYm7NqKE0h
GMprXEwW20HTIPUS5poIRjtc/NxX+PLkqroC2JU6frIMY2wpmZlGI/ESYSLth4YZ
3MB/dHdnS2Ia7w/9fl9qU92K+/WsRmxw8F6Utjov0WFDnfo4YKmWTCFLYTqXVK1E
Fjq+fLx+ZWsuUEe//DSpTFjZyi5OgSrvM2THBBWtnMvd6gaIpDkoNnWYl0XaPKlh
WcJARVGvdzc1Ns0ErmRFykdlUtQ/mzKPmZY2nOVczBW8ClpvM2JWqFJ7FMlzNdlw
OfEflt87Cx9AV8F/XUncQf+rP+eo3WVVW7FR9bBBrqbi9MNC0jC+L5meaWcFh3GG
Ipvcm/KPts1MJrlsibwzX1m59BAZ9i+6fL9bCXDlYZ6ZtJNuuQPw06yz5AkjPxMe
d7jG386mRxdc8uFrtUK3WL3KNabqkZDvyoRW1SDCDYIHbfOvyALtMMhicYZtHGzC
RTvErV4BO7sDryu+Y5IijUKDidU9eCZRbz/vVKpmx3PIMTdg3R4tSUOzNpcnGv3i
QfTuuwfQ3WLQIk4iGYwNz47Wl9dkV2q4ICQboFeUAWn4Jaik5JsDqCPvb8Wm2jRt
WKT5Uo8eYPKlJFIAnjHvqZAJaYUhd8gwWPB56EZiiVdQ8jkEeFVJov90Kp2E1O4S
oAYRTDd0gKt6CWxxACGhFB/5o+CVuY7uZClAr13LNPvp37935UOZMrzVO94FJBIS
NcoRlHHnBQDyIU8u1mKV8QLuYWqvu/3QNCGekDRJlG3UqNwVhWD1QXIX5dQwvGW6
iIXcIF37Kwt6OpMwfQ8h1BBvMNfMuvIjUkrAVj1N9qVpZaK32KOm0NdBNYYcBTIv
/I9oaDQ+izw5fu2/iCB95IXLIKIXeVgm+WwrFKEaQdAB5MdV5m0aRlwYySr8Cf+S
Rze0CQDmdgEyA/JrvHraDwnX5H7r0qE2Min0BMn0l8xJH3aSlVkGEcJZZcwuYJl8
ZtAJHnmiYuGIqM8Y4FfnUqEL1C0+dGjkQ7Y6zVRhFK3y3NpBM3GichkAeUR5MAw4
6vLejVtYSx3q7YAyd7AU3t37bS9jgpbib49H7cwqQU6daDL/vegrq+TUUTDA4FIr
2XcFaTGg/h7RGzgVi/H0ZR1HZGJdtW+WqisGlikYvhh+EmyckTAoV6nTMDEz1oFF
RsLVoHWubcBGtHXfSOnxnSKGOzqsH8LAnnm7QT+G8KsYiDQ1tPtlELUb/UtkVr6G
Sa6mMc3Ts1cTwWg2P1bBX0FRqjbqC0netcF8IItyvalwba/2LWoJj8hN6gcODMyg
3XjY5Ur4dzgVa+S9Qzrsz4FLi/DYxCcb8taEHbj0NZxyhBL1AjmS9UVCNSc8uoCI
2HmemMsuo9xvxTFhoQ6s8tjIKFbBHXqixEy7RwcOmjqOpFLNq7kq7qmk7XCWKwHH
uaoYmjcuoBzYCYhZm7jigKqu/75WJIgQf7qlGqN0rbnxz92YC+hUIWxv4PA8fnNb
Mh8EgjCvQg/alb5jhW69I3r8u5/CpBR3UJSqvNxFjPViaY9p+81sdumCvvboGkoF
UweT3GfmvZ6xgblHjac4GFi7fPk17O6alnUsloeCa/L3eCN9/R192tc6m4piJF9U
6Qo2sm8EJbijjsDvfQB19/bW6LKLsm2wVXahklApzKAliawy+roYVtC+V+/8Lp3u
e2mCoiJJHGfAJpkdW5A0sUmYxh5e0uOgXfzPU5dXhGV/4GeEMZty9lIk8Kej8lgz
3/BNUpKDeb+CA2WUBlG2IiGAl56pP1P7goIU9be8vwj/MOQEsmH+E7tF1fjK8bZ8
PiphDL/EwiR4EFeR/BJfaILxcL1i9Z0jEtO81HNVTLyLZZHmq0p+G1pnQn3gUirG
Fxjnd9mzUQTyvh00sWknoMPb7gcRQvh8JcGy26q5TUUoOxOedlktaQtcTU/QdUrA
jpbvVBrJ8IpM9uZKi4lmuJBd/u+jKpcA2wc6nO/FGBYlhse8Q/AHL6Osg6VXIYdA
hY9qTPoBU18FGGuiGNVrNM1HqZzTJVkR4Wa2FGQGpg5MicfswT+eEKymDPrABsyO
htLa+dlOd5iNI0n1WX4xyBR8AEn9H6Nx6CF6Ik5fqYtNihcIGpt9KwfpgdINV+0S
RiGjGJQLY701nPSD69fz+noXnn1RdiYKThqRDb5t7vlCxu50VV369tZTqS0RTgST
C0IWmBBZMWpV0mMiqPnDEoWMxFYgZLdYzOKQOxxdazZWIcAXqiAQexp7uBnJ+Oa6
B2cXuxgKQsGaoBv9k1FrRjLDx4M7z8IMiCGcEjbYLgagB5Hi26BlI4suU6+No4AD
j0wHLcvjLZ+uhJJd59eRzWvAQZt2oEp2BpdwGchm84ovptDuAgQKx3qDajmeEVpr
jJ3ytWqH3ZlMj9vdHW7wNYhWrHUt7PC/gOB7tVj7nScsVQGFCAevuubqYmG7OMM2
EraRasz0t3eVmBnCvyipxTbmfQ62HPBJMvKlwt+OtlSeOuXU2Z6X04Q6w9adjWwg
bgGrkNEZs7jdnfppoXBPk7mwinNYGtoWL8bnfe/RikBg0kG2gH2ONL5AsKYGLggz
5dyH85kD84brhGc1tpkEHqBSBAwr/HmLluGef1lPGgXsjC64xJ41AW2sSIC13Ran
Up9fAZTl94HRLoj/MbO789qq/+4ofuJzxEOCV8hkcB3eArgVcpdPSCQgmTNPXjqX
GPa+pxJpqbdxxKiMIPCFH+8j0jwcaZHXJtLx8RRR2MLIVL734dOUQBk1hUgyyCuw
rb57na+RcyazkA0G4FDVv6gsC41wMV1F7fTfh8eI3Xc+XSAZn1bZWQs6osFKtsnZ
GxJYBR1u8ZBeAbOBODJi/xQWRkNnC5xpdKMfJBXxnwwGzINJgYrD10cNwlIaZm5q
diSl4jrbcxrNi/L5J6NVPAEtwrStVDGF2uCKCmRo+HV202KN+cvBHvx1e2N0mPq4
RkUmYiwyD+8VwQAB1MwbZ9ojsWQIuRB2VMjeLWoijwTWtLkmI2tRSSBS24SEfLoE
e34Ohs25doYOb36iwAzmu0eIGsjuQmcvp0KGRc9dB+W+8mibUZepWh1MerUYGZ++
oXpkForW7o46CcQja8lVw3oQRhwNPVxUAMm8nFw9TsFU0Ugwy6ZJKu0EeWTks5Ku
SCdqmSI9IuSJGBPCBcK1bPKppGxSUj8xRM+63MIoJwDOg7K+H96iNN/ZqZ22Foxl
siwT6/ZMMgj22Jggd9950+phnC0zynKnL4N38gSjlDKdsHfBLNYuucOrBQ6sS3Dc
GIiZiHUi0YOsTdlIsvAt3TIP04YmoH5Xvnr0Q2WT/XIN+GCqk0Mz1Xu3Xyq8Dbv1
ljQpeJJ72HyGnE8P3F44x+7hdV5SMJB60o6BIF6PVapgvylEHCmcfeAmP3qzeKxm
9Yp2GDCkrZwqhX2Wgg/Akn3YSyIbFb6TDlwdrXvHPpBx9M/w3lnOOyJe4awU+Vly
eZYkTkL9yn1P5WL+ZKLE96V1dGMo6KPyY1kiVQ1+JdBF9oapX3g618sePEixnB7J
UHhkHuDsr33rkaacJBbK7e8V2Cv68kTULpGDAg4mCLENL37UcplHoVkLCCqDUb0g
hQn4a1d4OWc1dB7vxt8hg+pipN1pSO/meqTlxMDeK2DP5undzHFWMoBPF4ZuuzD3
Ny5IynI0BL6mh6cqBNBwXSuRXPaoia4BWPySCDy3VxKtCEQbTG2Fcs9+2EMfVJF3
IV0pmx85oxz6MVJxl3Ld/qCrujnRYP+KPKh6+sAbBAqATwu3WmLygDIszMTJw6vx
fb5+rZhcb7B8xgmt8bGgbtywCq1fZUzmWL03pBLA6MG92YmphEYexBhwDSscgrwl
Lqfw+4uzQAYfMAMFQRIQi0g1vdHDARSBNLGtnqcitcDq/WyNyu3PuFvuGOZpgJgQ
DGZY017LMxHpPOYo20Ud6LiQse4oUkJiuOjMQekdVbUrjIAaMZWVrVijVHvodAcu
CntoQDpdpQjuB6bQUqyRocw0CmSUbHkLZM/vuIXumFrhdKVswMZlTrXevoaIfaUC
0s9ooBrCXAdXbfMWmdOc3VBXxWITK0cOpcVzAiaQZxjpfixD8hHJQdygOskwEF7x
JH8uzLIFfeGuaHFv7tDM5VbpQQLueOsTn159EiXSS6WBNzcE4Hy72EehI2cCc0F6
KmNoNheE2eM8E22aMcMJ+Eg5eXwQnBnZFNhu/S8pZzlXzh6yAPULtGMWjh9iZq4/
IMDPK4b7HxfE7lJSuj7pWrVOd6EP91t5/5XOoa0xaZ21sRpgIYnd02UmGuaVZemh
AUcX7WXrcFCVFdF+wp9A2toBMh1m1ZMbyoBWonTWqNFWYaiwHPAuPQxNFl/3Wxp4
4fo1xT5im4PZZPNTPBjkk4Y9HrdBMPIFnrQaEJsp1ZATWrMon30e6PcSV7JB1Ot2
7s/hkSK59ic/XJekiAwgpQ/Xdw1z5a1gO1q6bVod78c1wq2gYtSIovPmrjSlnSQe
APDB/7OdZT/fmJQLw/RvQl4t92qlxKB9KTTbH1Y/MtBj9/w0e07ksuzsAdPKuxhR
2xapJgK+1jfOnt+Y0v7ZALlc9pBg0jdT0J8eKLfis3jYi2dRyj4z40IkGzur67Gg
2SiZIruVXbmyqvXePTflI4Fam09IM29u9Ql8OihLKK+koradhWK0XBTKUboodGry
DxLRdm4UZWc4/x1nhsGRVzlP0vQUphkK1ozbdcX2/heMT9hUv471z3teWb1KARcW
IeybJ/S1GDDQon4n9vHRGmf0GLmjh1ozOe4U6SEpHMINP2eKhNHk6PF8xygyQbpE
B1U0CswjK6CP7+x5Yh8gkEiba253aSTSRoJs/hchW3OfGqHvwJqWigB8Bxpm3wwj
BgG2hIojzOQTHHbjZp6utko2UsrKLCTJ23NzDN+hLc1jr2ICQssitMxaJO3cxn5F
xzCYmdfVlg4GeGCYCyERgMkUNJ3rSHtA+dh4jUqZlOqE3kZxNBjX8RoitQyU6XI1
zWiQ9Wbi+l0a65JAreciAe1FSiOzK4G9hpNnQola7dmN9DizYHk39kOtgZb3TXci
BZ4jOq87UWSh1kKwCw47a8DKe92lhfN+yG1MWjg3mEwwzMqhQYfkTby+xF7PE6Ct
OiAIzZy9NY/jp6RiOaSel4lJCYZl61XKKOx8oQspvNgol4IMY5Rga6XrwOn4Cfw6
6vLan9DkJSQ86eejWcw5ea2x9OD9NNUOjNcnwyrmBemZv4pj3tgd6HjNtc21/pQA
EXJdkooLw6nFhkx9Zms5gs0R4FNzoXiagg8KSVlxuZ6X6Wb2Surw/x9RpiohFMCI
DtP3TSkoP10/vQxZRz7esTTS6wFTL+dGX+9hlQsxYjhSOzJtZ9d6/cewVspijZrG
7nSkiHqEstwhB03jC2IDhIA0/JVOqpyXTKSwzQzC7E8Fu9Q6mDsSTRXhkc9961bQ
YzNe0J5j2rkKuj1kXw9PVRZCh2SGpB/zyAlwFRlXy7gMTkMQQot122XWFhEM/NUB
r5bePmFhVu1cz1kK32uIBDZBvIHYNZ9TRQvbeBXHE8/cgbMkw273rSnGt9UYa2a0
kGLG9A2Prpny6q33HHsLlM6XtfHoPSdLvysGpt9ELK8TyqVK390OQLhODTmhpAOQ
th02670W4JBOmTJDJieLucgDW8TS0RiOAGUIPDNw9PW3FgtsYrwj6TSOgQhe3unV
7r2Gz4XuicWA9aTlRxMJVQR+qwm0G20f5IE4yxNr1SYYQfygReVl+q7ITmTt9lzw
2vpQQA/mSgxJpenaR6Ze0NNhxQU8zniF2htR2EKhMTqbKweBcLWWGb/qvtmv33ts
g5337nBmsKhvcbzAcSPtmsdkemBYMHoh7e0FPdZd2C9C9vzZ3yRMfcRz9bQlVku5
Gn5e4pn0/2mc0sHqLIKa+QDXVwigb87fMDME5SFB/rCxG2tbXjjCBRA45ZWHsBGv
lenpOOSmHwxQbd/QbyMwVHcGey014hjlXR2jcjeDPG9iY53RzlOe9DmxDLlgjXYC
xhVQ7sicZWa3bmoLoFQU0hBDg5rFrQDjQPnorel4bPQY6Hp6qLgCDJAogLX3h/37
rWRrlZou0IVL8itET/nnknowNbyD7ZcRz5VG9XzUSQ03UXjhGHmczmp5BMh1fTQX
1B0rgOTeUve8sVop80P6SV6MaKDZnD5gTJQoZx1ULwqTt8R+DyVHLnAI+9sz5zC2
JRKnLy45tGcCumiyExz+Kt7olqcePZ9ik889xVOatEwcBcVYvuJYuMlvMhGdbzYj
5qGtPmMITLtiBPk8NK+aZNIem/k1NN2YJFXRjZ8l1CvfUOnDZe1s5JSa8H0nfvqg
hNZWBrtkPEHei6ZSBKl6DjfKcKKgnIjFit9RismFE1BIKrwS3wsr6jqRzhS4ebRt
9JscHJhAi2R6bi9YcoQu1ozErWkEQ8HATHes5A9FJ23n3rtFDBCt4bK+RFTjd1kH
z3182hcN+H+SKJ0zX+gQcbaDTThR/87smQ2yWM5s4Pbp9kDrD7M14KirQT04NVGi
ZzWI0txnR2jfVFdV3dlsBkLm78L5nZKZQfFqeWUozEfq91VXCF55Cef0OzCiWy3h
jkp4JdxeAscxIvuaH0NteRKM9fenmr0M2O3fPEPw1ZLyRnVvVa8PnFDquSHOWyGy
8g+voUlGo6IN7wGRwLHIi7b0t72tKnOmOMYasweZRcrGokkokXEucpSijkUo+L0L
28dSiK4Sun4wNSP0tdomaqnE+zNce2JnxY8aU6waQdu8nQ19TR6lpRgkV4j9p5Wf
58bK+Iz6sUG9pvMrB+/YAnMvSAD+O5WRcIysBlXObPQgG5/xVTcCt7Zm/Xa2LKgF
HExxhM27Yk0tffhjIiKbBl2zH/qtMJA+VZxRzxnFN6a/hhUhiIhcc8WmOGkPD+hf
G5bQ51omuCAAuGuGPZPUoXNm/jGjjlum+9VF18bSEE9T19OrR3G8AwXWmILc65AW
Z2pEhPDM8fyzkUDdoBGTI5ED9KW9TqqRSliFfersRDrvQgxc6tVR9ian93qVYpOk
knJBKCIGQyqWNURvdlp7hnpOWsW/rvbYNfN3qPpp7jfPE984nB+2U8kPVtPpL7in
oHtO8L78PEyur0Oe+mhcicwd0IYFMASrYfc6SG8h5jcqLtDnNFJhbnP3A12jWZYd
5WyHZ5bR51E06rIHCcbSBCDjlji+q2QcgjEea9C99+WHIDMe+/PInJB/9V/TVsJc
BHOLbwu7LNOX6Iw0vwXcQqrH/fd9fwo7NnkDfOblCfAFU47uZ7IIUe7gn3ixHxQ1
0y6m83A00OPPWGdy59LkuDAlmnQEefCqv6CqsFUjloSXT4khenYgFssJdaXkGDdb
1LRXvM/piLNXb1giSkZXDC7rGdPRSLeWG/aq2pA/xGgq3ZvdehYFp5OG0LHB3c6U
FWLHapUiB5N3uW76xAcHzwLDA2HonC+Sb+mwXSVkNp8wmrb1VK4YozUNNH54pdca
puFq/wN6/whKOFMu/9Jd8uZzvpxwFzUFWs+RWpiW0YVlbyxxRNnKaZBDax5H2Xmc
9R7aoJAN7GyOHFxvnrbikrhIe37Dvm0TkbQw0d7JMBr3Wa5PmqDpl+SIZyIalsQs
mUYPivO8ZEmD3062rVsDPbVTLSFsu4d+yLIWjF4gzz6YjPFNNUeW4tiIb6X8r8AT
/soQQkkRpdsXMwR5EO62mqB7+J/LTNReVLj7AJU8AT+K263VHAwriPIQyZj38Ks+
pgaeHP40TM13LByMYDPzwhehEoyU0M63p/FIkD8BAFuUJzRDxG0TP0jwGaOlYHxb
7aNKpoD26rRbF4mXWX2mysvTe+DhWsKE612/Ut563C545YpOVJtC8mJYEscMJTIk
17BG6EdykxO5GXcWmNpRSlYW+/v87AkRhScmpB8ntUCgTxibrQIXaQSwYdY4S/0b
MA/iJsCNh5u/2yUE37t96AIfq660sscs4R3kjCIPsZppouLMBRI7MYAJJalPU84m
60HuOxfH1S3uX3VVqx640SLR7ZP8VB6VGAL62XV22K9uUPu6We5BNDGXJANjaAja
QR5WNPn576eg0eGUuItlKYGjQhXILigOJeGDtpm0dyWPR32iSl9T5OMaIr+h98X9
IgaomfzOPMCyou0dAUoy3FNrywQ0c6ji4qtJoHIC7GZrswGPQ7RvgPG3cjr62kmO
NVBAzd+XRVQW4/893cIMjIEvsP7SnmrtuokvslxOC2OFKF3m3OvZANZaYysptwZZ
GVLBEU6VDCIlDarHKtdN7VnKAiTthOtOrG/8qhD/IaYUWwmjgE/RdVq7/1R1+Yk4
fXJH/poqmDcFlvH86RCANzcY7hw/GYRAiayZP3RKdy7bUXOA0yOy8FuG7NEGS4V8
2Vij/U9SH++w1G2hA17dUGHNdSYm5UKc9E6VKDl7tMnyQfXirn/wxhnLnAV3HH5C
dyUZ3cznP8lGmfo3cgu5M5vH3FFy/eD7IKGgj4uaS3w5KGf7U0pTfCNFRsG9j7Fz
dO7XA6uGgPjIN3tdOLzi2kXTiwiFkN5BqtbkMma31rICNYz21WKX7PwmaA3Rm0wo
hx/SOpQJ8fSWqVgrpTAdS0M+5rlY7hWtzk2iHlO/Go6LigyZmsYfk/w3S9Mqg/Oc
GPdzEBI5eSKD2SBKGLWCDa7gK4TodrquODcm3X+yPxmXjiDQLFYlTPHs7ZfDA0mC
8p941Qm2obyc3WGcV8NhnxYyYhTIPR4VZzJYp7gLTufdo7oGFYzILYf54Bvcb8lZ
EWiCNCesrzQx4MEhthqWObAQ8bHAWvLq63Z1WpjW9na46KnKlpo9S6Leb1jlcGRr
piVjbsqPHQTw45g6eL18+pI6N/pu1ehlVBZXkfeSpiVp/+y5+I6VZru1V6J53gcW
IDDrtENyjdBiM5fecNl/HVhXYi+Lctqn0/AB5v0reVllIO2TlhMISVZ5ijNZ1xvj
quAu2uT/tAobup6i9qU+P9zjsSTLm+ZbNqQ2lg3q1urw9y2XRkuHPdshxYQbkNh1
b4ho5WfsQl9C9Ra54RCTsto7UBiO1Mv820+cVQqE/HnkngfqaTOUS1cfnJzeO/+s
aeOUabPTPb/NKJX3uu3Subn5UwgN2YZ9UkCbKxI/cQW2z1wG9qANzQfmejINQ1eM
GJnXEroxvUwyfO7xue5uKVEREnwyB3XckR4y5aUc8l0irt4XfEiODtowvIOS2Op/
XvUO5j3zZDRn2mZT3LLicphXLBIK5f6yIUHVnFamP3M9GrPEYOXWM6opNh+LomaS
UWKAtfZtWujBCM+B01eMpLxeGzXIc1g70wxnvW7a+dtYrnCr/fckJNLs7sfpn5Yc
jgGGKPXc7MIfKqxQd68cGvqGVsTsyQ4srSW4m/Lsne9x4yE+9r6Y7++YSLVcFJO+
rReMgFIz2TTABdaqdkhTRmPDnpK+JaAgXF5mwYb0tEZ4KScwWxOQZeZEVUAuzYBk
Y20ZykpZdddPUQ4502+j5dER48Lvs+2gAI/zkUws07rt8rJgjHJXOn/jq2eaO7Cj
WbuyD+jF6eNlIj+F5sEgmdwCHOc/cATarPkdCNuouh69zlzsmL36YpDwd7+jlEQi
uX0wDyW9P8pmS7QfxIqQLVpZu/lxYksJDL+bSbqd4Ky4BO1VSuzd3iDZmpxy7zeM
gZdhpzN3NJ3SOUyiVXX7H3WyC/AMWmpEW2Er/6hsFjvUlZAWPl1DRDlq/EbSu+O1
o5viB+RzzIWwIOWpz6U2VLy9d70xixYkBTNknAtqzZpUp+4mPYgQvpBDVPBu2Piq
+rSDFDEZk+xDrNgcTEXIExcowb7E0ar84eEVmontrzemB7H5GzMIvPAYm3qQrVik
w0O0SWZxwm2h9gDDbXQe1MSGBvqURHzWVAQPjI8MhooZZ2ehzaIxPle9i6BvFnWx
9RfK3lsYwdbblWagY1rSYibmYze5J2BafFgdQa1m+raeXbh+Mfuu/SFgn2BzFsNz
1HaEonb5cJxaUvNM+mksJXmUsaHOcxRLZuAMenLjGcUabbr2roIh8QH0pqIuAKw3
/2ym+toIplDvT/tl6RrX19EOoZqMiwf2htIEA7o0YC1FJ0pYEH+4ymIOy6BVYlkm
PpAJH8YyBd3YUDBbpLH3qxhu0DYqDw1jph5ggd5ogcA/fISJGiMShuvm3yUsJyEj
TF0xCJUirPHDHcNFJdrGOzyvxTKzSw6u5PizQbAHdB6TI5VCUN6ZNT+RiqSCWxIC
tdVD3ysDJNX4bVVR+Har9qtZCdkiu5D+4vDCONuIrGvxCaK6jFc2s053UhOphsRG
nQNHlVIwJscKnAlVg7HwIsMauIMNG6l06WUzSfgOiasJMNxkIif7grbLQL/Wy36k
zWqea8YJPnEPLHGRlchT1H4oqgUpHIjZ+T+jbHGhJHf4ixxMmC5/Qb04nlr8JKLb
Dhgo4orZe+a8mKM+cr1qcUlEz4TiOwJAG/yKIL+xTgAgVSJpowow1hOQYqaH/HS4
rloWGGXn8oE5NkD4FeA0CgvYrNQ0Jaboj8XbyGIbHPUqS8fFawF8CXK90xkgItkX
bqs0W+RAYrqrokm4QWCUojJ4KZKmn70aMdBVsMftcr8ljx8kd4nnhzMqFmFmvmEW
aBB2d4goNJzdOfjqvU3IqciD4BQwt2d+3DAbDeDYX9lBJTNLLCDw71BC3qdhp3u+
KdM1YVHw9kMy5G75EvquZEKy68mLNP4rDLl4PYdyyPVccIBNK1D897Kb3sv3harX
C6RmfGSuqdieHIgmjQP4JSxyOsSplVjweYQVbkHDb3nbM0Mf1tb4Atwor+7UER/R
b0N8d41WFh1pgSzE1T8IDGti4fPTRoFAg7lgEJBp8a4XAoWH91IkuvCobEhuX3b6
kcVyigd1IszufGQhS/pWD+NhQ56FrlnQRTdgcAJtUvGjXNYu8MRCwtR5ZU1Rx7D1
KoaCKLQMLkQm+iP01+VwuRuHZmm++oAUTUsZ3fgzk/UcoIcXX2tCIxSFlvUlFUAp
VVjY8+YoBLIayz5tJZv/KMoOYf4XE3qoHtrR8wCIbCiAcyRhr8ORFdJq+LeWvN2Q
1StQ0tWyMj44Gv4LKkow9NuMiQYAfxzXvDS7SvkeF7DnF4A9U3xBVEbRseUZ+gFY
Z++copdM/D0X2bDf8zFqC3jPUk3gQBYpRfC9eOJAaaPa7LeE+KwGSqrJm2Y9e1wJ
WcYViJVyQk03rnnv4+EmfNGfAKrYt2MUWuE6Cj/jDprQvYBvWEipxo8RDGd9GcnL
NTD/yaUnsBCQ6aDCzI8L+WVGaz3Ov5hkQBrn1bG027sc5Ey8QIP+cdTzrn8Vr5VN
WzTij2A4w34RElCQDUjQAJXdKmO2OJE00/5EH5+SpJW/kbihge/ltMVKGfU3FCUw
z+NDI1JxYszWxS3hc36pCALy6YzCJJVDJC1WjnyY21ctXYgtZQfdurKDpMf4Jtra
KIclGmEVxnQ+3j0thIgL6rtGd474SboI6usp4GHRgsPoYnIsPPT99bTm0JqNWdXI
N/vB96Troxa/kWIvGyC9sAaYKRT+QgMhUBVROJJGuDZTj5H18I8F77zBWUz86O9v
FbxnGVzJskPki4mbCGA4HoDQx+BvPgaqvG51j442SNvFZo2IVYs7WQOmOP53PoZp
jS+R9pkL/w0HwdpLxxAPA4Ah2YM5P11fk9K7mypkk0hq1aKCfUbptPuKFTb/F6TZ
2QMGiOhEgxjmrKcYr6mJ+C1ZmJ9cx7tB9wlNzKyowmaYZ9IF2jQWkU66jHPzvmHh
ViNfp8SgtiMhkJEEIZ/XV55Aghx+VaNa2wDDQFXzMitbVaLcODQ2OjkV9DL9mSaC
XNwLLnS/DsvUDn5bZMg+/6nDE3Kw5JPP8wuPcw0SYfSOHSJBJg4Po2us7QoMTbAE
agIePVSb1LeYb+GFD72QWtR3Q4kN11MIk9sFWFqHyVF0XzDUpZPs/aOvjGVAGt3O
kDhtX/KWwobpOmtN5MJ5oQzE3pW519rOu3hNsNquLDlcLRtvlVglg/WQUTKqIjvI
FtbtdrKRKjhE5BphGLF9J0fTN1eNcOYVVu1tWaXLnd2pwHYEb++o7fIPjaAa0T4K
ksuRVwAShGVqcr7f8cR5mMU+MXpyGfu6NSqqgtidqRZKYXkPbpJrSYvGCK628bNz
3k177JaGWeU7mnRoPC08g7hUH4KjhTEiFtfdaccYOt4uKi34uM9uEpm7WbjlvIqk
VJ+Krj/HrKIdmromtqdxy0rYy7ece2ij5hcSL/P+cOcr1U26k0WYRlOQ/nsHtglL
o2ALvUmyaIWJo81F+t4pjPNLwxvrP2kfBtaLKfztnk/0mNU9vjup4uqwxSwy51/l
/boalfqiY9JeL/N0aWMnjxyT3Yc6+aSIrIJA+hfd+DZjNQ46lDJVEU+O3HVRIHR+
MqCzGhRN+KetibwjqgCSx8+SGuukmrk0Hk7UEE0r2otR7Gu7d/mD91eqA3V7PALY
51Gpixf2/Qe7u/zX1ZVDMNcB9nJbAEeK6wjJIcO16wvZMz8tzNp9cMAeeOsvZS9s
2bpAeX81//A8+thMkgWkE7w/MuzVbAnTFW8ONaMzNaUFsdG98JiKtG8JtOCLd2DQ
Wi3oGwawY1xK/TS2EcMMkk0m7j4e/oZunHZvA/OJO51wcgPx1dp1MTi5ChJfT1Ld
XujG082nNO+7GORLHTfMUze9glNZb9dgXWE5SQb/Y4owJPs1DNr/S5DhZ2kyWxzB
oIyTujSLSAkSINTylTHq+8wWPbWx79WwnmbHRhIR+1XxsHeyt1Bg4XCxHsbkkWXj
W24+R57zwAqNYNAeV3EW3j/sIyImkmyuwpZ6dp7NO7NJaUbaVc4m72bocxMuFFEd
GT0kL66uS/ofU9US+zsO/6peyFBT8URQkszE+gxB7ojs62zJriHamB0xrFuO31LT
ifYv0upddza+LpHzdBpDPUEFnL2VFET+ovvdXcXiE6aAJMcvjM68Sfd9o1Zx/kUu
DkkRoxrvFwWUUSvxDyGF6wbbfPAbEtIYuCFsaP+uHJ4gVVks8j01bDo7Liy5vBfr
4Oq1Ts5JMDJISg2f5vm+sVVQ4ONHbUx8grw93tzvRU9laor4CMGNWt9xsXIIGpQd
PJGWbdAIWn7PkBcdSnJ32vWjYYpgVyuk05kJlnVeVkudhtmNkQxR16JT99pbsU7C
sSpbZC2QB2j5+3nQCTv3+v+FXTeyMICKCtXsg7YeB0qJFpeKPVbtOiv3BsD2yhSZ
1HPHG73HWtJjxY7tjG8hEM/NKWelqpGnMXYRYYNBBpsLAPHsaUWFMlPzKOXvP34j
5S4jwnD9uLgyFKrz46blSXIxc9YdquZu3y3XOITvgq4h1RQztw10bJIBzO3hP9Is
xaJUKIDC+njRs40VPTMAUX6SOj4uQevI29E5Z+ubfDBOLDsV7iD+nVbfW7zSD/YF
PbBM4FvpYPBdP7Nl9tnmL9/7bGvzyzt4/Al4hkSlRIEzRzZYJKIRlGcHc4S23c85
YZoTNr2ll3rsVMg+2ijtKRtjRYOOYLFf0nwxL5aj8yiNeomu2Qm5rDUZeIig+2z8
97cErlJAYvtdn9ZYqVC7P/hUDiFVtDIGLf0fb3AzevwnwIVPi6iUXnYuJcdZoEvB
CWaR75XWz2g1sgGYU5nLEYDflZ2sTdfF9DvNd/zfwRhUcKH7yGfvzOmTCLyDWJ1f
mMXkBJIJCsQ6JEwhBq2JG8A+2vueYiKFcn5djN4odZwOiMxsucRpBFDh99LjrSch
4dvdkXBtdrd5waMsHyurIPiENiBfkTDBZR/UZEKiNEQs1ONaYUHm0aO1HNQIm068
b8VNyAqFgRVURBEXBvNq+UiEH9+qIZLl/MDMvovpSWteoCqKsGlEg/+NcZ7Cj3X1
TIOM1jrSzf7+5cL2MWRts37+eD9hGuVfLBwha8RljcGEwFfxrgHpPkTkDWuLDGHN
OuVoXShdd6gwmGc6dVruY1QIvtZG+sAG8fpLtg+OZc4yJqtAfQVB0Hdq7jgf3ljZ
BigLsc7UB8erqoHccusdt9m3Pmb9Fmd4ZOWRGsbGuiAqmK3iXYC1MSIlvT6ckEzK
YbXHb8DSurj76FBWrSrr+/YQ4Qks+zQYljVfX/0CIhYhhLuwRMENzs04BRZCRpI3
56eGvQftYJM/8kqSzmrHwF2c6SBic2PeVY1SZ+F/L1J03am44yRDlJTVMOvD/ziJ
SVQDrJ+YVcdHfbHIam9jqH/taKVhLXgybLhK5UZC6jZHUWEv4jmSSgVHC92Vnc0c
oSyJj5EtxWmvtZZCBpoTKmSY0qqWJup3VZB7+f3uKMgu6aKsRgkO5qd5Wk1+LFiA
W6MkCgKET5iLwBvatUlH+CgC6SCltwTp+CqnLUuxCyy8wMhLV1nXqK6Yv9lzCWO8
D5Q1zKfp5mk+euwrZuUK3MBXKzPWgWbszThgfkPh+s5fJ9B0kkOCWrpa4ObFKz4Y
J2oWxJWHTAABX9EUv9rNhMUS9JNrKkGj4m06S5owdawurr7inf2nijUFUQKwEAuZ
/me5Ch3mKHDOS9eGTxbqfQ9ufkIvJGMTgblLzUfVwy9BCd3ZHgib6qNXV2rnBv4r
Si/bIOMESDFJ5kvBORB0qyysATgcZsRkZ7qaBJilrDsa2R5Ay6k9HAgOWFoDlhPr
swWpTd70V1jNXkc+8rJmElPD7CQdqRtqLcS+OMNUiLE3OWEoX7obufLzQ3GnMRDM
56PkRhn4AHLFavo62rdNyPakY/F7HqhkRq2sMmfMuCINxmqExB0IrvkYG7yP52vX
k+FvA7/6jfzoj6G3zI9iklYTwcMJ8GqGaKS9xHOl8ghpq0vaJFF1gLTwYEKG5J2b
eTe47UdFA4OzKGGG1jxgZ1MygBMzz6kgsXPbMaDjyQt934HgX6w0dDVAMCroAzJi
0duytGj/IEPrf0eGe7PZonjw/n2nIdai+SWdBgG7GyXOsWhsHbJmUCv97lgsqSaI
M6O0lyJW9vwTXOh9qtwJA9osxfRnW7NwBp1LV3gEqaehy35nRLRtzxy3B3JAFRgv
1CKtDEnwYkLcD64r1mreC+pQQWZZMsYgncemIudHrSBfG4Kwzw9Uc+v0h4VqVXis
FGw3xHhBrTsXJOVK7zDI7JTCnbu60E49OTXZC3Zvzv3IwIATorxKlSiutaFJJGFm
6R1XA9g0XHGA/+kKYSUFL+kzdfg2EJTHyxT6BThJFmjDwKno9lCp95nW17rcJLX1
NW+gp2E/Dp/PJnaAAny4zh0Xtyh8eipZV9uT2Ptt2wGA9GDxkHTm5C045YzoUX3Q
rbP7YsZJC8ADA2fMSP+ZB4j30WJX/19VamZ98S60RCOu20Xh5G7thgyH+mhOifiR
WqpLUNqQeBAbSPmYPgLObqCY9v+SsN8WgarAoCpoIgrMMeuNdoSTUhsY2nozbY7q
3ziaYRfxKhiHnzkwFbz6m6NYAiTUSReRawg78IIO4GDDIsFPD0+ciaSsr8ZB1omK
RrZq8cBMje66Obl46GvXn2j6pj92lx8Y3m481i5itq7hEdj+8sf6Q3qIW6B50YrA
OKqnthAxcwO2i5S0XzWUFwiG6FNre8WKKDkTuhNG1u8Kpq6ERTCgAr7+FbWsreKb
pKdXFN8bwOB1pq64u3dYL+wpqGWVmwW/n+CSwpIgXZd/X4s+vMeeXlglG+CJXku3
PDBOEzTBKo+QGr2zRYPVoNOBJMZtDMQfGtDGiQuJgLqZnSurRYayPGtGG+tWoRF5
Xleflo+7eLRfSPHLKswZFukOFRbH0fRY9KMAwWosz6LQbvPRsvtIvfnxjKaqUNmU
NpI8Rc5XaPOJfMuKXvQBVEwOdzJayuqpQ12BvYIVauVTAwzO5wFm3+6ZuMH3E3E6
1AcDzhyoaHVg5HpmhR5fP8bKbTxH2nTNLig5gl+L/9N3FTeUTThM46zJH5eeBxSB
b+ac3oWT3ABbkQ9F7C5rO5iEY8XzGi/ZW9JKdNIw9RHYVk4DMBnBfyGF9h/rN2cv
rDe359N1wqrPjGwJXcahf0B/Cp9+n0K4V9/IGKIB0LbCeEYvI11Gcc60s15gPBQ4
LWDA5/vsogC85kudKrYrDuk+l48n/cmTwkGUBD+u8/yywpJV5MgHSeEzJ/84C8ai
cwC5t9WtQbPh+VbgHdjdv0eCiefYk25JUsve79VavzdbjZwT7wiMDpF3m7wfKNKp
h+MBtDPH6I4TvHbA2jbqxLBY8r5OEOLjjsAp0teJM23v+WyWN1EOYrP7sOl858HG
PCO+OOGatRi3I5RjFfpXqv0iEWbOcjOt2I+0O93RdCsOOI5cRjOO+gjbStiL6sIU
1YXJC7eY/UeJfC2r/8t+4uaVYt5NRER6zY/poocK/r8Z+8h8Otq4cp8ua4u5zvuf
HR6RXIUXjusdhkSIK0o4I0nN9xktWKfxq6s/M6db1E/hOTiNMrIoxVbg4M313x10
AHgijmx6qo6PCGgDA6pRPDf8d2y2kjxLtWhp/D8EWgvgNWRkDpdB7ottw3Uj9ALK
0PPjcsTHn1qC+WJw+sZHdVWzgdHOPJy1d62vmWDOT+OHW5vZA4rR6QYG9EXBFky3
bpankwPdVvS4U2b9DWwOl8giEh6Gt++9JIGU+4LAOYastGQGEui/D72OpKFnXY6W
Qd7Kx+1IaClD0G+n5DKaewSmhO6Op1c5Ya9Obzxn4E3d3t+8CGfOtmoKhXTs1QVu
n1XzA1Ss3FKuPkeLaPdtIRhY3cDbVq1XnqvwXPjDR4Kdjw+kTINSwrNrR3I/YzAJ
8D6TM4hukY3OSJwfZB3omqVSxjqp1hkSwcjaQ9yN6D9xMDgxZXLpw59wbSROE/09
Dqj9zOJJCXwN3kbsj65q31IdmTRiY8gjcQtdbfqGiXMTfB9GYVRYHBwiGmzI0C6M
D6sYBXMqEzetzDfss4TJirDrFMepu2kJl0vMcDo/E4mJY8Rj4qe0CRfWE6iRAEKS
eCwjNae9wX6z7I1y0mX3xwYFQBXxY+6MmTevn0eOifDWfI4YyVEQlxwdjk4gpBGT
H+RZLojynRiKBQegpWWRg1jIETSq/lgSBnK9J2Iz2bTwd4TeB+9ccNWN8B1cICvy
TCUJHe5gBXgLYy0mx8MsuriFPNz2zpCG3iBJj3IxCDsoomlhFET1zLUip+S1JLKB
fyYgb/Djj+a6dsHMS0V1DELPTpUGNiBlHzTQdkb5AoQpb6OE/Ym1YyyU1PczUjXd
iR7+NdqYke1rIrbaeU0+EEZFC9oWOmAbhHOUB+eTWoCLsVvFHen2a822dQlPKyR8
dP5o4rHoa5CUwuD/GR+CGRz6aKHiKxzPGN0BCpPzpF8wro3odl3tA0OSL4dPjF84
0MgCNAaMsyPtPrjvpk31c3/JR7JapLbb7ePwj5nY8EhmkbKgfyGuPn90D784l+4m
zU7WbjXnkFOpUAr5xMZ/63lG3bahqHwjyuwY5OfpCueK7X4HgtGdAkqxgEYr6PMR
T52/8CuQwX4rTrHVGCYGQxRHduGICppwTsnmvbomZ3f70LveI42ECxARQB6bi3iV
QmBiDNPhuwgXqEqlIgRdXUPo2yCLDOdoj0P3OIaMMW8kEW543RGu+kHjvSV7wlog
AnBVwY2I/SrB73XE7wSktdTmGd8VD5AUbgRaOBY80bnKF/PZL/5Y8388UU5U63zf
BgzIqZEFmgX5UthfrejyaKP7RLGvjofhVdJlaPJ21ovoBydb5q28sxcuY3T/pfDt
22TVSIlV0QyeiYaWbJ8s03QuRLbpdjyLDJMZsF9mUmQ/e7dtRLKQUA0btV5xJ2Id
UCpfSZ2Jdhh3hFrRSnuI5Vhg2aO+ZZweW+OfFtkpFO/RqBh2VU3paoovIAOFPuJZ
6BoP4wbKIOjNhKwAjO1JC/1qL7pBara5D4S7wXBGhkVjKhHmIZqqzxv2psZw9l/E
Y2xDDroM+xiHMP3dAmjY3QP1NEMs0kh/V7a0Aj9ZaSAm8t81zrdtPl1quztrNw7i
vTzKwdO164zWn2RK9pG4jzSmgYjk5YgEGiPF2UkYjeEbuIr0KeDO7ForGevg0aLZ
i+aQOe4wV0aKatoLdujI1Lswfl/RkJlSTGcrpftm41IAQOOY4cLdcjRHMpoZZIkj
IvwJWlgJnA0XUqYncpc6aHtM+QJYqzUwoBmmatVOQAnvHEJ4NgVaCr44HoRApKWU
8LtB/CjR5W/slYElKGY5We7kP7g1IJalGZkr8GBm4vtgjoXgFqcwcEkb4wUB3jrc
eW255QXI717DrfMe5GpAwe7tc7Y1WtSfypX8FxJsHtD3TXB48x5A2qnoikqORjZA
TKi336+kULYWrgExCW0LjbmFza0s55JBL+Tbq9UnE4NbQIUXj7qjeEJ8kSHQofNA
2/sLBRzVJanJbLKu4otw9Uh0TK34qMEzQu2emIoEpoh+g0EXkWqrOO1IGHW/myw/
myBKmte7+La6gYCTnsCE4d8weB32SW2GD0x9H+cXJnULkmIPaMuCXXrbI1C6KWFZ
R7xcW2aKKaiLeznzpFIjTVOas9bGyCGH2kIZO/WrhNOjNcLPgMyVMm7YwZF9PoYi
SyXPTnpr6C547Hz7k+AZtdtCKwfd0yZnQPugg+b3qSijQhA50DFz4i9O1ZCF8Td2
YAwecv/g2qJ3ncmtQw80w4P3Zpa0PO0j1hZf/hb3jJKiG+hsbKlhEI9dr675BGPH
lsXhvv4OdGYVjLtJ3V9EjZ+4INwsFALJVRagv4vnd8LydIefZj+uUHcymAsmcq1F
2jCk7vp+/jcPf2SqoiqF/zyi5I3GMd04jhGQAIAfwlAk3mumr8Qr0HCsD1zQ+3QJ
L2okJSKWO4pJv4THptYwHrr8pdZ9bdaUacLxb7Dax9rY7evlh/MRG35zf5Aafh2a
NQvOXp0fqqf9H0rNIXdpMIRTA6DzcVlpLQgjCuMzM7wGW494Eo2jiRmbvJ8ZET0M
nXj1CkILvfNf6xO0ibn4H8D6jKoue37zdEwaJkDW97RpDghRUYOuXoTKlqaQiQlp
jV29zc3kVu8Tk6qjBW4O4l9oCZOMGaQ+Ml4AQW5VtH0FXlVOzFyxrGjSnD5719hJ
xUEznZx9BbfUFfWB9RFwI/CznP7fedUvSZomvPLwF+jCSOZo2nxKWLuHEfbNhEfy
VUOqmGupoD53NK1d0pOlu/ZHNxyeKnZCD/DynKPjkyyNbyMF7eCqenV/jx+S3d59
K03uK+cmg2nV6klykVNp1wCl9rIndcjln1AKpyyULwRZ9c+or+kbT4cQbuQpNpnT
kkl37sy0oip7xpdV+E0AnKeQQTiNduTQSPXC7yaikKbd4AFVDdYfvE3J75vgDt9A
DH/PNzdFUO8iybJkPMeIMoUV4a+ghqQrswW1H24x7b5Rp+iyx/F702lRgBPLPK2x
FH0gJ5oVepbvXVYOUcgNGjFA5F7joITbfklvJ4A2/RiElsmAVjHNWMVTZ6aRHXcs
00OUtW3PRFJq7RJYU4PGK3XQIaf6HxymCY+tri+v7wbuoVrScvhgEQKy/w1Jly/Q
K1GPKbNITSPCoufTpclGojyn1OjcKhOyPPiK5uvhj1HmiGu8U7oOTmY1eqd1VTAd
Imj5FXwlS55Pms2KlwV2pt7jByhztvpbvuY9IxJMZntB0Xpmwz39QULApU9J2Mae
3ykFyMQ5DefTuOENMMsN+Ad3OCpyUWRvh+CXGtW/N3OvNObbi1E265ZmmMm/pa7o
SEaV+1opYOwk/9LwB9MoJ7oniWQe0uCu6VVgGFFjJx4R4/tb/kW5qwDb3ZCEb4YF
Tjl7L35SvCJqyOrMpxEGZEbwYjvGHKULq5Kov4Gff9HyrFitK82msZI6AEchU2TD
gVNPnLQRFNXfvdu0dwF7OMAyVPUfQvtenq+EtBJUevsY6NDcV8N40W3DswQJvtVr
qO6hrf1st3+dPAt0w13+iUclH3tUfHjcHvmT5A1OPN9JAB5sl+mL15o+1Z26+2C3
A9yufAoWoBfJATHbZwyfKmOef5kbAfBxwrdSvUiyHUOso/fNP7UIKpgnLkvzWQMa
n5Z7lVGFhQmYi2QN1Hma4hUWPg7KvJ+UAum+xOAWGaYWZiFFt8gyrpY0fPtvT+FP
45Y650Yeb6aOoTaOLVoDfmo6KJ3FsL+aIu87O/wVbrSV3Gsqyo5OMPdQmeGH9LCh
8gWq5PM4Vi5ixhSIY03DNqXF7MDl5RpWLHn56Pn8eNzA5od95ow9pGfV/NZRu41d
srVuEp06P+6mzfLcuKmcbXDnGx+SQsP1rlohe/eIQs8kD4P3Rmjk6ZhMgcOGaQ2B
R2LzLk3xv6DJlW4HUhUg26avL0FmALx4Sp3hS9LJxX2+xVdss6kdK/IgTyiY0rLP
KTw6xnm5N6nqBD5i6kD3LK0IVG0P1GgJj7dxkFDqT9EQsw+UG3qXnx7M5NgzdWXW
+AYR9+qJH1HO2kupnQRyaJlE8/CJPdnOn1vtpxnryQmPb5NLzM/EY3omFTCFE/ni
q+3ekQxoV5xecD+DZ6ecXhLd6pqJlK1DrnETI79WZgxl42YmP96mUNNYIE4Z1gB/
KseT0xy9/RLsI0zBPev99cCg41JUk31aqSLW0nXw6EgxbceFtJ1Q8piEvFtVfttx
zgeWxhUIngVDqjH7nLXQMDhk3y2dC+MqIrlnx24dqNEfqZFRGcq9+5+pyZz9LBBy
gBCG4x90wO0yV31fmfy0dywl/MZsAvmgAgsrWUY49D8soILYAp4kO7Mhq/g9z3Nt
xEZX0ah5QvxJD3ip6A4/GWY4K48kAi9gepbDS2J8qnlVss60CAKjTj9Lkrtk+uDZ
NBmktgv1m63yjBxFA+g+E/C1lo6y4WA3qb4JP+nMpr+dzDMNqJiIs3hLBFAcBVPP
a7Q9jw73jHRHS+WzY/tv0G6spEe5adsaIctAq1ifMQR+GfsYOBlFPTjgSg0axHM0
r3CZsU3FPGj7m8d+dU1qbhhjoTqtXjfg8ziIBIZLzRQZKaDQDcf+OyhuoOulwt6y
nlJYeXtuxMbw0w0p7W0/unXpkebHgZ8W+nRanAXidUKfd7BJKWsFzqpu5k+GM3aY
mMXNPo16zfP7xlQlYlckUrnUbLc9DZEqI4r5b4+EfOO6t6LMeaVwBhIc441stYLX
QoKfMp4aD+aVE0WZ23z0I3Ppa2VfOEYV8mg43755q1PMXZxuGMJYUe+wGz7Z5kY3
DuFPOok/r+A4c9k2dJI6l3EXsmKNv6KrGk8kjigKGZPlSRzARmFhIONQ0+wGfGBU
ChzFn6xbCEWBeM9TiDogSXMiw91ol8/N8QG1/Jdr64qOQsWHeE5zUuHkXrwgvula
/e8tZ3QkZ9Ek/+DwgbzPI/d1zelPBLaXtipmirib3VwkxgEhY7GdHvAqXz+v5Z84
bTuheADjlYL6etoYTxbWqLi9p6ZnK7tNfDzigciPM1PqUrkMROL0gIYGCttw0bPP
8oxOR+1/Bs9xSWAo2K9BDcVNl7gar1ei4C7S9ushC/OBA2kVTPFr6wO5eYf211XC
1hL0/63mxL4K+y3KIyY0sNHU15mrcIqyXEAyGO+ukA4HbIIAAvbZteeCgch68ZKs
jvGHYUq+xKQorTtROQ9Ln5NJGZUtttF9YCl2B119gBwBO2BJtbZAjkKDHkFHXJWR
S6N1IK1qaajJfoHzOMqrlvGe7RCDGiakcnyNw2qaZKTPEXXxbm8fZ92QAgZIC0aM
yPRcpYYF4QBcv3rcWl+O3joNbkcCJh+yKp3GlaG+mIOij0IVwCp5xVQLlgbs4guV
zFr3xhDyNJBqqQaHr0TY5Ks7d7kfbJ+WHKFOIXO/rizstKEbZOvsqLkVKtiYz1JI
RCv3mh427ZtefPIsb1lFHRjKgqMuAyFVt0B08we/kxZKhcAR3Y6fBzK5Bh42nsI/
oUbmk6ONH+C8rZVf4T3MqKTgIhSrod6jU7f/1FSN7cSBeqcrOOb8JIsrze2mc6OJ
fYKj5If5O7MO1g7p3p9fyaVrx/MdXBR0kvmKTkX91jzE0dSetPVpjAiTjdUEldwk
rUDgaqSw7gnwqtRXaywxsEqZlF32Q1TiF4Iqar1qf7Pyz/P/WLe+n+15wFEluOcx
smNPAkUOtvc3XbzhGrWL3Gqua5uiLeX4hFtHXoE2v6Y1vjWglAXwbC8VGskALHV0
9k3JikVUsC0kjlwc7202T7iBWODBbt/PTxNsmvs4AS62jH8j3OJ2d2edZXYS8uSs
3TtId1auBuDT32JKSaVSghdRZx7E/OAiG5usSCHrAyw1dBXO8dcjMpN4shBvRKEr
LeKUJzSh6FpHphCHlXDjYxUcLOuDjbzifhZ3WNMhSKYmD/1PhvudEZWWscKj1OpU
rFg8or7WvlOC4kPkv5feJJ2w84rOo3EdwMImyddmGODVmCoN66f2oDc5mxuIWnBp
+Xgf93dw/O3CiJaMErGj37mjG3sb+lqetX2vgs7qgVHXjA6v5CcRUOMez9sxHBV/
2fLrdSAoRbbzkCzWXyw7YtC4UL298OSv0zCACkSEkgepSNUUzBpTmea+0TmMIWqh
ilOVaeDvhsGijNF8M/NeDl+KhUDinDgEYM0+v/IqxTtWkWTq+Y5gzZDLv+aRIcvp
rnWLeEQpDBWBgR8kmq0v+0EcfFQdZ8VY8B9jQCHd1pPYF+bS2gDUOXfdQaSP5mF1
kqvAgq2/L4rQk47UD9jOyGc0Ma8FB6WnpjuqW2u2Ggz4gzQeT9oWfCDZ57XkAE6d
5vsGBZoe8v0SG7nTloi05yQBM8NrIlPTL5onaJFg83OrUSEhSfNLdOOE/jSbFOe1
eXcKJmKiJ//84/S+goXsJPSWaKYyhIYETzAfLyIov33cQr7RISzehdBwDtSakmnq
Cj/TybWj7dJX1OW34mi37Zin3/xqdhM9JI3bEGeLnltb1uHU5o0PpMg4WzpqET28
rrDQKFWyvMF/N4R6gEP5tDOP6qZHqXHqCvO0svKgfwf3ecIEFAnuWD7xHrnY0+wo
evmI8snV/k/+2523BVHcHQvUwJJnYakMRqKPuuZlXoeSl5gNSisMV3GTNldeu0Wb
cKNrkQL1aMQVQ8oXklI1Rab6hpbXYjea1G/mfLuS1SN6g88twmupM03i5eb7Aloa
z1n6f94eAYuVKyaPC78BXKpRmdzLUA2qwfUTfxE5rujmAF/34tVhy1+6qtIAYfNl
opbpIojatZN+nXYmn3P9n5Q7JV8DNiAcSz7ASIvzOshcnMPqO1we6pf0copKDLmE
vyIYe7NRGT4iFXD6msYmfVkUM7834jQC3c1AX71m2A/0LlQDmzeKd/DC4FTuMa5k
VmmYLslj+2o/e/jzEi6lOdpLq1x+pcPjzqW5uc81uaQei2VKBEAIFq3ejbk2sDnf
/edaJy/gHCMMwwQjSFwrtnlhvK0TKwt63/V8Yfut95EYbS3NDpPyj95TIsaAZV+H
DpcKGDn8qCNHV4nOV+uPHrjkHe0oB4y5DEP7OgNwyW/wZxqWdXXvxG7bT3XRnpsQ
e+ZGKftxWJtckHSloc0mQjB2wkjAOwSvJ94iAHUD8FdlD0IsW071CVszPmIh3/lH
YrPS8F94bLA5XRk4SxrzEaSzF6ossTAquvlBkUyuhucbjDRt3LPq40F9Po0NxADB
RpMAK0k3b/C2q6acvhbOKKxi0uEG8vmSkTt1/a5pIvh5O9CAFNLMPtkdyjIlBHUO
e1yTokzsO+7yprMwdbMcnZTjP3p+Y6u/4acrHRsdR0QRzokMe6gWyFLTlj81rRBP
i+lYr/gvdxeokUM+yIipaBR6SUcVpRVKsRYLP0G8F4Jq8Ukl3WXHUDY0BncpzVKO
5SJBTekb61SUqK4AhldYRxbIJ33LnqRT2FGsVy4wn0lYrBfN3SuhKgZ+vWrg0wLQ
N4r00FQR16YqGQoF//LVyBHkYMXolH7QTDt054/zFW0d+6GSM28EAuF7iiQAEwa4
aGMESNxjtnuZtamVXcznqCiIer7F/v1PnDOc+ky1VP4uZie0+ReM7U24OIPLOiGU
MF1+zUII0/t4TBCW66Uhw/1hdD9Qt9m1Z5VY8fz6hp2cANr1LkfVP9/Vd9KBTVTm
UBD+R5Ao9whS/UBlajfUEI4JaeLtIUxrfD93emFr2JBusLy1yIlzCufsODpcLKir
6jU8PxkL90ZuxcmeqBgKOaGYxwp86pC12Ke28WTFM4voZAr5hng9mYnpk22bvfco
UiZ+7muW4fi3QKnmFOIx73+01hFQ5MTSAyPYl3686DXXA26ZTT0aaDE9HTgIblVz
v/nYXXUQT+jz3VgLbJBLTFXWDXrsy215YP0ETP8GcEHPalumB00DjD7iYCSqCO+6
nhEso7sllrp5PnJsZJW00mwC1ZhCkWD/oUeI2W3xmyWkxDZgcMR9Arq1byLCyLr2
uRMTBjrCXIBeWsaJuOEbcaSytDH8FmVhFmKA+DNn3YpPJTHXRwf0khNuJiwWJQRZ
ym2bAJzMOqiNZjHDjqGRxqDpYzkEkBRlOwVdHvSGfjFOK/0u29fDqthghhacyzzp
S8/dZGIcpCwyNwHCp8LPBozqqTJpS1jkPtF7yizj1A3cr9hTWEJhZVO37DUrU/J9
wqJxwdmkr0UdmZanBDd0hXpba1KzQ584chq40zlJHEJXCGtCUfoaq37dwPL+MYpw
DANrOI7HFBQQ4QkGWlTcOA7JxOd4zvHhKAGutfzZVEeqTbfveAar+V12wHhg3tG9
eRhvG8BmZ8LlV48iyNxZSeVpv6/aAD+iws1GdeCoA2/nJ3HwgQBb7IqBcmpErkok
qNattkCNUmHp4+NHoIr/gKTLcsRiS9sJJB9OE66kU1sv6DtkTcVgw9kbAic1me5S
mwASiZ0kNy+Lnc86Gs5xKdXDQduzy/R/Z2SdDQFZIiKqwe0RysCwuR71DdMcy3BR
MP9S1SNQc1jXgo5kOfnJZoQZNj83CemJviTbpB2mY1/5RVQUpFb79XrgjjHupZhs
eGYuweePNURXboNI0jmdW5dHHuOY9sQDC0+CMbpjtu8SW6pcbE4QeuNsfKAwL5mz
qjpj7mJ7Yjzk6h1DJmijDbSijtqLthDsUruyUw18smrD2ZkfSQtpZ193f9JZ6/f7
3UWXBUqSjX87W71Zni8RfLjbWIzAET99c7kAqqu85xmT5OzMrzbYoNsBu7i7owBc
eaLgnT6jCXZ73zY+UGKKeM/kY+pA3XGCedQghLYuwnWQTUM5QgqZ1uZ5hdQoSE8n
08JAowc1hbjAAamawNgg5zNxHVMOQiKMRBuatBo+whly8XRrbZBgSEgLbqPi6TqD
4xyXXeqHcvFLqIBm3UzlUuUtrhc51kAjWCpyw8H72Bn8o4RyihJWBi86YIeVHtAC
y7Fgve9p+8cPWEOBEglUElLB2iSuQcJqMqQl3yJAQHsAoF+Fjv9FwnpkTQs1uptw
oH5xi6yYARjcMYbOa4spgzkSl4j3BuPCs6BuJ2JehGUk+Z4JBvOjb3XA2xlkOjr+
vI75ePey1JndBG2afCKVER0Ej1S/RsmKAaEq+ak5u4m/unQOyXfPs9zPzdBKl+S+
GtVyczHh0qVLRo4jnaWCmRnBTYrbbIBtqvKFWNLPZc+LS0OhDKacrsaIzwW1wNg2
/WiSkWQXAXgxIGQ19+op8AV+b3WE2vr19lykfO8c0ghGUPY6alytAjYV8mH4ERzv
/1AMpSTyRZre8Uxo0a9AfOen7BgWc2Wr7VbW3e+A1NMb/WjYMxXbtW39wMkqiNRd
buSqPG0dqTjnRix4KQF+Y/czOTpCWFgRx8QoDrKXhuwg8E+alIMZ76GivLhOpNB3
jiqsOrF+WsTwoZcRmT4bEViw33rKnLax+lww3GVJkOU3pos/6Zb+FsAy+DJI4TC2
L4tbmw3+qSNfQ3yhoLtVdwxuELGl7nnzHAU+LhVRCDv1B+3cOhMz5tZB5RseRJzM
FnFfC1nvvbkuoTnpbaerQqzRUKmF+bFCgOopQFjGmmGmVylKWPlihsEdxhRbqaR5
Rt2qMKQcxZs6Txrb8fs3x1u7Evd49NbtGJKtnxpZbVsuvNK7clUTcU78R70N2nli
bg4K8TTgpGiy2orixJPIZeQ9CwfNKf9TRqlQx0Mo6kjR8IxAUWtU3VMH1jxx25wS
ICIaCchzsl4VPMSdbKkI6UoiPKe0/cVVL/q/3fM6noLtBZCItimujAkvhNESgpIl
iwi2NyaCFBemBhaz85x41HYi456Xsg8zOhm468aO23anQTLccSkwdos+Jy+hhvmV
Z6ApNuX5bO/3u9OZww7ux4D3799xG53oV5F1q4BFvxs2gKqVHhXDmxgxChP5om4I
YFhxTdXxCkxLaOpzUANxRWKht2ecmS/mhL3jfR+qMPjkRcqsVrca2ksikleNb268
xZtwYOpBwBD6W/O7a0JJynEU6/2lApbLIazFDqOi/ELqW7j4gzUoUrCriDLxpPPA
3D9uQ/d+ZD1th916aBHIfu/b8pokHehVofErF2h8GHyrBa/YzTfLSRURtLEuMx9m
EAcXLvbamLEqLtG5jl/B9yUvjTfRtDq9W74XHYDEJXkrADlehHmAUW4r/WiMr6Xt
bI5a9+VbXBQFnoCh3d89jxAqmOcMaacXVvv2KnTWAEfSECooVdpbgfKing9ue+VZ
MEEWkEyOyHWavVq6An7ysOcQU5Pz8mRrblZBMg82DzWTZkeSnYYYQ5LqOgnYhJu+
JVEhgjpnriLzu3uVsiSLD2fOFCZw+ACSdML7Ca+hWvNZqPAvW949DmrCYkkwV9q2
sLgjnYz+A1yfnucQEGjyzn6BOM9Dm2c0zFWa1q34SuZxkemK3bUdGOSDoqFhfMeB
1ZO1qex9U6lI3stCdbfZMvs/jP7/TYDSFF3aLb5JhF81OBjvGVLN9Sws3IuW9ybG
Nx7H6Ujza7qHxoltJwpl6+u+q7hqLM9TyIdpytJl9bYMypnD7SwOAfPa9Cv1xYos
5c9XX1PFLyzGzL6ajO6Frpfgxk+uILZiSw0wta7c4Xw4C9xtOuE/5ZFC0z8V3U5z
dXkPO9zchWlQnb/IKPDR299Ezo3QtLvk2aJe0D9PG+Y3Wu/8c6LtZDWoKKQ9vB58
lpeIGFbmyv0MSd81ozIvKlB87S2xdMPI+7RqllLmY7I3MkReaDi3oHYsk0sD2+2r
3bWdVc6w0vCFhySEOgHp6VIFEOxMLyTTXk2q6d6bpXry/XCTKz3b5Usn89iAFYfR
IsUopWzFmMrcmp4zcfDBCi3XKNBoJb+GzV0q+AgGVcUxJOmTyoifW6YyNmnCTEXe
9Kp/0Mc1mHY22Re6Kkpo3DPM0i6XpHW72irjEYEoTfhReQe/pDYznpvVXTqeClyI
FTU20BaqYL7sDypCMNlQ89CQYjxELfdN+PjwVLvU/lDoVrYACjq/gIDj/AGZ8ikl
5ir0aqPpwlOGr0d0hTKsuF5Ae24aOXujSx0i49jSYw3DmEjHVeYrih/lGOIEUi0z
hTtuhQyiFcwneWi2flT3TcuEoLC1DKznjOjTc8Kr/0rVhgCx/Gl6cWF9KygGyKyT
05U+CNku5gJ6AnwNt+XM2YhdskWiO2WbTXbCDbnaSk8Bj72HdxT+TTKlApKDNwi2
Y4F6iLwcxyLR+fQcIMV7p4e+biXWaruQKtu7z1I0W9nAigiA2bBNoKldfZP2nyoJ
Fs+s141Xjdi2ZwAqBCYGdZ1pxRCQcxGOwd3X0ECJQwOlFR5vDMYf9rALlhyRRBPT
tbav8r5hCGm+5W7NW0btE3SPCHQZRtcb4cQuCf9RyniC+coQGUmH+Ps1sj1764cB
raaV0XpB4ClLQVBEvrn+/gbcPmPVmLxuX8Nb3dpybNiFR/Et7ICQFYJv2Sa7spNz
4S+i6YbZmZdRUI1IQpKZsFh0X7kfFzTKKv4Xp2aEog2VNBgS8hxDdlFVOrxHwddA
eUftt/u1G1EiEy+IC9QYB7uauraEtnJIANKHjaVcwrXk/12GVJrElPTGQNTp4jwm
MMs5epmb+Y4FF9I4e99Ax/bp9tAh51RLrULJduskCkRBhgsHIFb92mDxoL6yiip2
34ewYsZfJ4H3ikN3ImSOv+tD3jwQ2cI0mPQmhtvgm+VwkWrPnVw4NzkvUzXBRWb/
16w7CozpzicEEJHCBA3snrRwu2Ki5ZWnxqofdoMe1hV9THaWSierhskRI0AlRA3Q
/MXn1IEwgEx/fFi8KwJKuUXoGYG6i1jjtIk+QiIWyQR3iAT1etjRm+ZZFLZSqtGL
Stj53HPVa5/TUaDeINNj/yUYoYtXc8+QI+ui7cCsw+osv8HgHBIUtZ8TQHjrE7rE
RZ1ZInPcKv7nCbpOomofTjURsK1NslkHzQG8tSNYw7SBLQNBGGxbnSqe3SCRTbOK
z3p1UV4CXwJqeAj6m0qX/Z/pGAjWFIJt+2qRk+vbv5duX25E6EISP5TFrZHz030d
RzLhvFQfdOgmHqxZyx9s+zO6jEYknRtEsSeoEjFYKXTH3nSmjdi/oWAFwm2yX8h9
pWjhmKrv9LX4HAXbj/h2EX0C/DSf3MTEyrtr7didRgjMsMD+pHpRMIKdvzr1PBQ3
ve7MVglYKLILnOzXe9bz2RpTfgXJiBFhPrMFwYwjkbA0Gtw+YKfsUk7ZUPQuVM6/
a3TtItA5FwUVujtyrSo36oPVIf7Xx9a7zhZbIhXJXCbDoip8hqIwIY3DgM4c7R/A
fNX7z5+swxC8SrKoWf7s0Tv44HvjKBBX8LfOhiM0hwE/ZsQ3C41CjyjZEF5424BZ
jP4M/klBNQ+oHH1UZLKMTspZxT2T9YguE4zCfLQdgsa8mHm64WpQjOMEJZsiJ4dy
T1H/Xt+mrg+G1HVeXS5WtqBGlL8axzqmr1o742K+VHp+nk4LkZWTiBQ0dF2DlAgp
3pvw9Abykihucaf2AW83mN1rPtHKWRL1Ve3ZnHO49/qaEcD8LcSNbxJ8GhedlVGr
eTF4EJW7vwTkc6mbT8rh8rG5ydMh+stE+xGxScBFzNSPM5TY/bLtwYLvxhEtEo9T
ah9LlDTg/izCq3jaQhFh1fMshjbpOjsb600jm0B5/QQiFecGKn+Hk/9UWLsw3DBp
1smE1s5IfE0PHuZ1wzlrko6q8M6maBJUw8bTYPp+p+SUrATyu1oaidIcnywCVb/x
zRVF4KcbTxHRVfWQ3qFJ+1d8DK7EP2+69XRTWQWdYJg+md0vEocmFN3L+VVST9Ub
14Qv+KnCk33exbHFQ4xvfn83UAP5cBs2JAUB0w1UUFNNq1yrGGfkfEyl3FPVCuYQ
f9/OQJTdj4M/Dr2QF7ut8sWFS43/nk6I+NL4XEJm6ceB07Zs3QdFwokmS/6UeP9V
oQHdlf/F7oXouPP8kgn6XqCsWGQ946NGnSDxjZ3Y6f2mtkZ5OmJ5hw5PVydU5jAE
Puym6mRWZc5QwhDKy+v9K8eamkShl0QeUefK2B4I/bEzUTdKPFMLU/BYVc+osjuR
RfzHoUoQgxswZntu4GGrHP8Z053/g3OTwPXxGmExnP10J3v4sJuAwC3XQrjfuq1T
KVkmtvlBBhheXdF+ebohTqJi4TYSMlsns3UPTJQ9L3RTjmoHui/GZ9SUghdTl1iy
yyW9FOyyNJRLY85v4H6xJWQLhWi4PaTu/RuBrRahIfpKRlyYUk1NivWUUnLT0iCM
cLHiorcl0p0PyxkGzcKxB6Gc7g7ffOmCmu2AfgL13A+A+xS5PL4VIh5TVsm/Mok7
8Ztx36evZ5urVssTzy9fCLBwpPIRntD4V8JwsqObu4KgeMQB9p21lEkpS6Sx8rQT
/oxhYbyp5/+AQ5INEEV/jWuAGSEhF/bHyRPu9jlgkb9MTJivAbDTdyggnV0oWc9r
agk3H6Y9eIreDb3Y5Qjzzmm/xM0Ifc8vUEadnw0/j+MqrbQCTr5Fz/n7UT415pnX
EF6EMHZQv2ZhnnI6kswWym4J+uLR0OlrCTngXXR56xsW4zF+Jj81hhTgpKsvup64
cDH7Fm2ZC+WpCY1TnutW31Vy50ZLX92Hk0GysFxU5HJwkcaot3CTJ450lfwQLr4R
XTZAOdPP1CRttfOwaVRF6GrpsAgPvvXe2V9rCbPofZ7F2lIjSmhDxqeENX/kBv7S
cVru85Uuk/6h84HYRzOr/tQAlZPdbRgLZD7CnZeKlMNJHt2NCmM90wwUg8RwJuFm
JcIgC3m0TjqH5TLJzVvCm7ePQs7/vQM9ZRlkxT1ZitxIKi81ICbiSkKsZkkTv3mj
n+Y2r98Q3AuzOQct7USVh2phe90UP8F9JAPAMNZ8OtzssRKS4Vyb4QnyZ/i3Esks
/pM0cQ6lwHL8p10n9SB4jTzsn8qPYblYthky6zoeJgO8TQ2HnGdFA8AvvlZHHFA4
oyGHK8xdBMabjoJnUFB/ig+moFcOI0J8cIk66CUtUXVyFblS3oWZYjsYVvJplVOg
NgLAPf1kQgQ4HHL6vvUbRsGOJ6U/O+fpko2LgkOtVuP1d7D+sw2JPFLSEmLHZOzG
DOMLDCK+CnUFlF8TgrWLCewjP+soeiVKMpxsLYl9oyj0N+41jTzuCD+ZHsBvOiZl
AlR0QOjNX1BmC3NATetsjMBZSXpkaeD32p/VQCvAJQbrLLEMge1ks3BW/z9La3G7
h2BTZ4jRy8kgj6iBhzp9mitqDKAB/X+R/FD6vEaZKE6fO2GIWrIVBudhcijv7hDE
4M1krgyEgSszVORbQZ+YDTl29TeDIXwIl3BAlENZ9pO3+xMrTgdoE1agtSkPw0wT
SQ+4E6jHlZRaK0iNgTzYEjUNvgm4ThrNmpJCe8MgZGsryvA95dWRXIY65o6DOYKH
yvT6WCzAX4aIZIh1HR7E1qT/Vbzrhkr3on0eRFFH60joHGTMgyIjsjWgTYL1zn98
WAnwb0q8OyZROwXcsdMw5HSrCTT5hGDH5LU6u4N0OeIphpnuEa53zkiCcjvtuuIo
OuTVI6/MPS6cHB9qVnOTOTPCmC9xTFmiBoJyQYzgvmSyAkOILgo0blb6CCqJU0em
jtXRVquiQJPDxPVWkPDGu0SIvGQeRqwdiJ1mWcigL1gvmRxoNjUOZJdP2dHmUfTt
spK2H1ikH1WO9XdxytNbAY0P0y6UXMHpRJphoW9bvPvSh9Jvtppfv8lerzquuFPZ
PFDv7EqryY0OdQ4D829YZzDpZAPNfR+Co53RmAn8LbOq3o7VZBkFtoOGr6OWGV8q
tzDo32ooUBFeBq2Miq6HS0Mg+ZI9nm7ExIb289T/qlkHm2mH+TfWXJvI+uZhBuKF
1xASG1z6A28U+3c6CePrSqZnFPrgTKNZz18iV1O9DRiCx8Q7M5LAb2rESxuUioc1
F1iASBjJrtQAe4HyxbTKIjFFyJW5m4YcL6b6K6DZFz2VcKnld6in8hTb+65SDdIq
isfhkzaVi0lWNhSE4A4hggej/1j3VxvBkVEBDP5PhO4JZiGbby90ij55HrhHY1MC
cStJi3uqmDQrm/CpM5jjojwDEloUwQkESq3kPKPZw1kAIO+OSM2+oVUIT0kJqIYp
/DrYP6zvV4nY2IqdNKgEV/EBSo7xnMMW543wybvgf/xeg4n9AEknptcVfpR86Xxz
+/REpG5tgoI0CHy/JsGuqM7HqF/92fbsHtuGiDIOaIYilPUCjlmyfmXVqsiejVMH
/Pf68U50dJPlQBZUPMlxTVutVm/QcZbx2oQiwT4zSj9Xi/VVUjuSKO4FseN1VSVz
TgFxPeTk1TfagbczLq+41j5olTeTh2d9qRI8gWAo2ZdhLqoo9PVmlb0AttajqhSZ
XxE9sC/NJflYqUAnrYP1mlraZqg4kJ/lJnnO9dLbosgmkFVH1WFz3lQM79ZsHIHS
sFH+F+zulUKESs1j12auXQa/1bPGKAD6go5IKuvrOpCcRZdJCrJQtqgYPb2pQOrm
B9MOLxAe0Vv1sG6c7odQDZDAMB1Y1aINHd/EIgV7xyjeBaqA3HCiGzpN+ca3ijlL
7wqVJpBKeIixic0488qdTYihfDYM1cFgauN2J4Zk8+xCezOK4aJ+LogVXby/HPjL
2bBc0pRq8MwWOBUdwWcycKk37a4GTIGZWVsdC+tlgGaWL8QRtpp+GSOoiJVIGjO3
IANYqEsTsqiAzZT4z/X6ZBVWDEc2sOBBfTITaGzUNqyO8PhA03NGu7Eq9+GVbfZV
7R0l/NsoX48nZIuSeKXH1/zP+ACoc71Qdf6opdT8tZNNvM0lkOafjHmzGpPIPYJ8
8pXbItSUPKos+2IlmZu2MVn6Y+qid90lBAlzJxqr2mT9Qu8YFamTunpsg82MFUEo
Vqer5wPA1xZWDc/5j6Vn+ungH+e0LG4OMFNa2wXILAlG2ChAtqm0borhGLo5HX2b
JR+XbasDoXANPpXFhwkfbsbs8tKVhT0YqVmHfyyXlJogq1pIbG86R2xl0sa/v8fo
n6UpajDBCEZasBXI5Ewh3dS4hO6GYWZufU/D8y9KvaHRXGDp2pptVEhruRwwfEno
6EIRIM5h53conQNVGrRWjfX1Ul+gOxO7ybCluJ+LxaKtT7Xl1XNY3kGRL+lWpyb8
ex3seGP7SA1U2OwPYOuMA1hoqkVlRBVYRBadC6boKM9yQATqMSKJyAEHRobc2xAn
a8DGnKTgWjFj/WmZ/OLMtQoKuvox+OlJUE6pE7j7d7qXAZKn92Rh96KNDCHPwtOo
qhj7bNVB533+RpodFs1XCiI29p55rtlqxH+X+zjugHIFcGQFtd1oTcjSIxRTf5TP
vB/u8jJmLNNcvfNP24+s8O6P4kmV0GIKM+/zwwny1EepLr2KSZbefMKi8GV/DL81
X1T7seHn9IORnCblsSxdME+rbSiAtt+MbrUDTpd8GceRdr1+jqlm826l6y+5OtoP
0NFMm7gxVgt067O3tBwr2EoDptcuHFtVxxgfyuJ07ViFwuZz54AR6LkPRysb3Hai
FcqgW7SOPcJ55TrdZd6K4R0m7rAjlxJKd1yYLlbH5WskqLG1w0xYWQ5xj+6/s4Jt
fv5MgM+T3js3qXdOavxHSMZ7ruhap451OutVQDAzf1XqgT118sSPt0WmgwWw/7Bb
R9LIiCEdndRHT5ePe0Kc7AMj0NV5axvo5+dvrADoxGC9pKm38m7v52fO2kmpIuPp
WOVICqjXgrWKTodYIzCZ2nI8+W3thq4xloScrTuU8e5O9ZMoEtCPTC7ugx/dZf9Z
PbdjE1+4odLgWhQI3dYEpLSw+qtjYYSyZmwM+2guQKdD2YFAhlmPCkUFAGiTLzjE
vsu2Nt19RRVCfvma/IC52REWB3w5H4kvn47PB6BE1fqnjq7DI0o+EmrukNuZPrm6
B4+W85UzDXo/W5q2lQisA+kCTV4Tfu1miiuB8xPKgbwTQ9VPY3bgj7O6iuSTnedb
Rk+01KUEocKGE81Io3oZYZsvTiaRW6Jmm6eJMzS5ZwdpAoq+xdi6FeFdSGEgRMhM
gSxOxcLn8YR/LTBJickY5bXlBb0BEUnstO+JhZUT6TH3E6fDc0Lm/dRxtgEH1J32
wBdeKRImA4uLEJ7SnjFzKzQmWNaC7e1JOoT5e84ulBzFt9Zrs4xYIz1Nq6jiW0m0
naq49fvxXgWfXyGggkm6yD0bCeHJZCsiJtitHki1M6eUDLk1aZ9s78+eku80vcvZ
z2nkEDQW8udSj2Uk9nWzEkMr7b9Hq9Le2iIuEYj6TUi2g4EY3ke6Cgs1npIPHPQZ
YuKWXt21+YSH0Iw3EoTTZeAHeXh2+EoB3k6WxYriI8yy7Hkgag1jT9TFt2rKDpFS
veKMFeAeqQ/9D3qlD3aJv8lzo7o8lgDMitBX1hgJv8pm8qfouaN7rwpZwTFt0z4V
O6zliKxD8HH2JBhZ3rd/hbpqUm2RI5QCzo+xmick88suh+dsv24Vk+Z46MEujaIV
ckFb21LwLyeOBrSb8gZnVCb5S9cqecatpScMmJXVnlcMYIj/AV7mifmiSxlS/92c
leJ2WVShjPy5lvDLtR/6G2vXNjwGOnZ6jwc2K8yTzBvGxCY/YyeQ5f1La4xckaiD
Qaqls9qTvGI1lfC/r+gwQZAjsEuidRMR15dM4rJA1rLTZTPCQdnYVcWzbK4TikXw
QHtRzOTcveiWEga+s7eeheARKw2XvNE8omEPLKkHoZuNSiOFXHKU7yJfJax6vgxJ
RkOPGinJzUd4r5y3bwhBGioXjnOCcIvrDNXH8w4oCSz0BoBp4FnjfMIw8qUW9H0u
NJwNrP816zjeonDnN2xlqKZp1GGQwwt3NNrLCjRbC34sKFGawFGZJAshzj0FKVTP
okQnkmJ9sPcVJ6EQGQWLrBfMpDZeGsACd55BIC2TYlGY7ug7OXKYVWX7pSz7OJsM
ASBus2KqC0rDNgWU0+SM8DmLz0naWCiMTfNofWaGrScNEqMdnXKtffJ/SJWqH30h
+c5gRSzGdofno7YXRYuNSz0L6McCLaSsZgYEUxHpuPRgA4XGS65BVEUN/8Unkhzt
JyEqnURb/rS/3uEufJYghP//aboCsrc/9scKiI0kEJJTBvlsDbL4aRVSO0Fee4xg
MgI1DNNlg0D1SuDxjNBF78kyLs9xxY9H5kvcgh2C15UZSO1U2PMGp7j/zqjjswtk
S6IHT4/Pw+YTxLgEpONWtiSKbv/XEP/EB7dxG+K3/gC/8aLk7oDJXywgIIzp4uL2
gK4cUo04nMrY/BYbyXV4MVgpv48LBLyCl+2m6K7yTamp7QWZaGrqDGZ0HsdI+TYy
05I5etXDLeG02lVUErY9W93QIQrLDAnvr6PH70tOT8HnJZJYrEFUBnOCJVggy/Ls
QeRrRHTcD6BJOzaS10ZTkShCzwl8x/F2vhqofnkDg0+p216ZSul0HmgCqJnnvgv5
UTC8IesNNH+ZVt80tBzIUKQnwaWTJmxbLLynuf2mr/pOmrJZC17Z9Lu8SFlPBmZ/
KAEllqSOAZeEvAyr9vz7u7LPtEaGhbVEo3B2hOYG22iXUu8+Zs8mSFJdujVxInUe
yP2/A7bAD5GSOak9a9QHGVGeVCEbgIzq8th0S6aB/MhWSMU5572kkx04GBvw02D7
TPJNr5kWg8OchyqNvn02hz4qJR0rCgTbxGmHy9KpOAso8ZF69ga52MvhCheb1apw
CuSlybWxzCgBHRAAz4QNVHPW0mgRAd+828OhYXrbWOpyxD83arsfxcuXy5U9OgSz
zRNMCP5Y+xtSjd+tk29I8+9MWSZ2QGNIPAvrk8gj6ECkdbNTctpqdzLJHc/Xc8DM
a1Xc+OwIW0bMoEwVWHfrxXlyCDwD69jyHuVLMdoAAFUwkzhUslT7SxNGe5HX3rr+
yepiE74a6445+ZEk94fDyk6xVi1NjII5McEWwdLRLBLluEInyX7dxpYjsKFP+G3o
fgihWvUs8xowF0lvh+J68zHqDkv8W5DB/DLlb3ZCkpcNOXGS+o9TzyngEPmMiNNU
EBa/tu6MOXC9vl/uPBZGOxNds5k/yAS8mrn+ENsRla8Yqp8I11Ie6S6lgw5lhsn/
wfEWFFPptyTPQS9wRwMO0h8sPZyJyAT9UqhV5cycdtizLb4vEknscCkatWw8wUM2
MNwc4GTDOPPAMtQSskiGdFYR626XmeWgpDrg97TAfGeOFONwom4QFEVezJeNfrjQ
u8KUVBKKQ9cBM8xpOnRZ0C4O9Mkx4jq6qDG81UxvFk85Y/skGAlOuHWR6GwIqnfa
xUsDOL7v249JGRa9LwhThrijwvFSHMdu2lPZl2ZRFhV6/WgNVV6NRcoTjv6E2Hn/
ukP66jyp0jVN6W1AffM6iSqqa+l32dO1e068R/FaSnDBXq5Jg8s+q/6ybSLDUcVx
i+EwPBosJSjHycb+ezYcQHTEr8EJTJPNGqPnh07R/vn0dSulEToLatOrDyHsSSLo
s2yx+arHfUZmndOzNrL58faDL0gm2w/LLWvvZ1ARMFsKcvZnumoebnkmeGOhjvwj
4gCJ7Swjr+ffcnG2viaeycVtZGDno0tGaKyFjLB1+AFJox+T81EoRwPbSLU70seR
uDZxZCKUpZVYEfGajq0lo81JQx5DpFLNgeJ661+fejW2o5tEB5BSGnzUu2gmqlov
TVNoJIdU2pfST7ltafbz3CMpbJH8mibG6TXT3+Dz8a7BdlhvYVYuHFGqNtL/h2vE
P4e7HIN4GNTgi+m/RXyHTaRwK83h9SBf2L6f46e2087xHUTKOgtRBwa4RJN41PwR
JSlKCw3I1UNvsUNFZTDowuJoQ/c/7ZT/7ICdoXop/cYPMXPG6deEqrOV/M3DadBl
b9122Lxfvu4PwOhpCz+qTwBM/73EfBDr+zWTFBkLQD67xHmRXfdl+/tuUdoKC5XD
sxwRp0JgwqhRiUsmlJW94qPsiZrM8xAAjN5ulFAq4BpN9NZ1Cka8aMctI9roCBjP
90G3O3jqYoqCthGChMKUjaVe9MDr+xRHfqjFGgzcxUXzjrHo4dTPLvW5flr1FEsd
/6FPkg8dlA9dF2uEgT1Feds2Ei0nzxQrm57w7y03XLwlwK3ke9vG/nead8htum4S
Y/WpgylWyVrb1+qXTkh0tKgx50JnpRBeCODcYS4xzWnr8RUcWa+QZ1bAhsaoOAMK
uyw7FHVhtoHJ/xcFF5UX95OeFFFRwXua3hYxSW6DTO+iNEiXf7DTCmzhIfIUZ+vw
YFv2iIKGVUYk3WfRh+/KYPPQ9sxlItcmROmTUmVeQogQtnGDd1pNjh2I/zQj6Gc0
b0MLWM7/u3+XcanXzd83JtmCiWyv+/Li7cUVuVBgNj5ZnO9HIDPPXDKTfgOLh08h
k0cob6o9R6XxrNET4zBQweYweWhA/zm26i8NFkVpH9qjiNNftNSUhD2fGK65LLyA
gTgkGXOEWmcsRygrIUqyunqKklYnOcriQOpVsNHYMajvWUjoWpk/qLFGOhGqRIZa
cLXDaOiP5Wg3Rhaub952xX0xi26fXoDxJbHw3shOk2dh9q8SQzehO6GG28F+lTcw
0j2g/LgoMbyAgMovwtpp/a+Ih+XHLBa27Onl90t+qdMx74ZvXWUd3Zp3LeAkESWn
kp9j3xthQTdF0TovTkgCToGziR9uiIx+NYZiNo95gOnty2KtE7s8jpYP9PkY9Cm2
1Nw2HD9sRsOioF7pnW2ZbjyVGABVxsipWedpWPJfIZt1YNM2k7DFhbCjjZRfo5E5
UyIwZC2rdmfwkiGvT7uQUULSriCggnvfNv/MIvtp4NjCAyy6TJtps/B2ze0RAVDo
OFY9hCGHzsoQwDzD+ukOurvsqDKMv6s1jHaXgeT8XTfbUQMZ/jmgVxfGXGGcY0P3
fPQ42TQ1xSObX4yRCsQC+CPlTeJpEBZmxbgDqBXsZWQdmcALirRUhAbjx/WZBj/9
nGJOhbfMwWC7FGxRtvr1s6DkZBwsKW0o20r44eZDrNjDY9FTeFUPgGnaO5n6YGy4
rQQ3j9zsClac+PIswVoIgaQzd3TYIX5YE4TofDgnd07445wQ3z+2XHFWN0BgWxnj
3oFyW5VfSfcP/8n/lc56VGnS8VskssQh7ET+WpU8cj9KKyPgpQdGkBYD3YuVjU4h
nU1+sc5NYCMabApqAM/hVOs1ywqVRsxdE/DyWWgI47MDCHif1rUJnNIdRhwrfG7b
Edqu+iCOgginmp5qZAWw8JvIyPcVGJsUy8Q6mGqNod3sTD7sABeHuAiK3kCZGr8Y
tzIiw+tuFxt4J+fsG/7wWs5jgzE+2fhi6z9tDDtzRibj5hpQ1wzYEyP+jZej6g+/
X5OEvERy/BZXpq1ctQM1OCn0A8eQa896vgYno3mz8n1iQJThHxYpiJ/ZpsDL3EPn
3/3NH3MISSAFtGTfEzhhtmiLYb2xiaYSKI+gHCh6pY+huJJth7SKgbxpoI5cUMvB
gNOUzjupn8bWRLfWabpwhOF8vnycMCziI/RbAEgNOcoLnpZOKabCGTfGZO2ODVdm
BjCBRoEu68WadeCECGr8YMGM3rllm5tld5KJakGaznHJ5D/eAWmVy7oBU11qG0Q2
W9WQB1Vmw1nxW+XI50T/ateIowpV8H22jiK+TyIDdb8x2rd7A6ndF2yALkBlOpDM
kbUWVygUTvp+UheKonYEarO/3ZfBJBFdKwB51aKgbErewhPX9REFisTaLVOozZFR
4R5YOUY0U+M8H38Fs94rFBYdoXkvWSxisBa6v4u5EmXi3l8fVlq9SkUKai/P3sJa
h+Lt7rSuF6CIqfFel5pEPBUgb/D8Sm+Uxb22IAeZV9dPsqFE0q55tJhZeiXPe3om
N2ywUnBp1gGjVfART1cS+NfKaX2Zs3Db33lixlaAapGVW91kY+kEOPN1XLBC3OFn
89Frs9J6tuptTTipH2rozK6Y2sFs/sRQrmLdBdqbMSxyDyLKadhAQ/HrPNbyV0fh
F2Y+ArejAfH4OUZszFdQiJhJAovf2hQ3L3KJHCUi2H/MLDERHZ+0nNTjmMAb3Emx
7wGfEkc+iNK41bsgEoUJI+GwwM9O/h16yAQnhmfXlOPCDHebrV1LdoPrc0E4ERlH
Ykd0IM0pqCMrSXyNgDDhyjAicXLBb8iGEevltr6GFxUPsKDGuAFePcrqjtJ7dgk4
Jl82si7TYxkf/TLXp9gvhFW71L1LhwdRvkAOcMYlLe8OD/BLfToP3XyCsN7CUCal
egKCNtC22oJdFnX9ER7A24oUxCjwMrPwroVNclgEK7LQnJnrjkYs9Sm34asNQIeX
jR3Nyeby+cUJezibiy4AssgppJInDKXIRBOYSuqUY2Nb1P4DQ3LvhsTIKGzJ+KBn
D58PZ1LBPmU2uqxllDYdiDBfZhc6DTdEX40xhssgjIRh20ru0c5aEWODcbbV49JS
9LS5Uu4ANUrzGpNWoN26Hi8keE2WI1Mm69uqgx4U0F5xO8B3mZKtTMlqdSKEJsLK
uUWBI3OAMiZN+08iZvnYfBaIhqQRLnWXfs/nKKl1ibc33KQrCJnIg7dG6c2N9AAw
BLxpiHsD3qd1xuUdnmPPjmsnH0Kfuacw2QjObXH0Fq97IcMnIKQgiqqgWEnQv4EY
mN4pAJ1B3omQF2LibcmSpqDOnFnJe1/kMcloEMojsII0EYKtXWD+sFP9RreB0jsZ
xSWFSkXRW3vcpc4DW6+RAwFPHNpAe8N49hgPFJm6kppZfKFHLScit9Is46XMHCn6
2/+l76K6znrsR4JzWJyk6Jol10dvAakapJJydT6q+ZasvYaHtVeynvRaLPIRu2Bv
xXZYs32Hob2sX+9vLXU9DnjtUKT066n0i202AvDt/IwKfPU8m+dHPnQh4uK53NXX
opfeS5ijOL4jkKaIzHfWRAFHUMwPwbfAc334Hv2ZJU129C17qXKXhsnTzh6UHNBz
34k7PiyTaeOXSBmEDz0PPQIYFOZc2m2ukN874YSBTWvBMgt6ZrGWWHcLvoToBAXF
04d85UzYEDQ37LZXl66/JdgYdxrkX6ADHASRDnB57/XsAqzyvpAzmYmCI2srJO8S
O9fDwLAwhzBiGTbKvw48RkAfqZrqjc3uJCHKQvxAB9nah2ST5JOljl9Ctmy6M5T0
oZzUFDG50TgnW0XMWwiwk2cvCmd6eXmjHF2Vqo5IKED7iWDNS+KLXMmXURndZhiL
gOiakp0hWtvKdbYdPDQK7qmlKxGg2h/jAvp9dncb8k3TPLQv4kvTnH3rGJ9Jy9Fo
Pj17j63o941O6cV4mF7sm487iAJYqfpACiaXJjIZDFTFRkJEqKiqvJW46bmIyYx9
Iix5TvYqCogBMg2wTs9By0jCagMbP7ma6/sebYC8v5DKzEPADFBg2tfO016gnOVY
NNf8fr2sJ8yyxj5wxA9+Gblh/qlnnRo/QwBl21NU5XroJ0ADaeL4Gzu8FI9+6F4l
pFLX4pDUsVSW7p+ZisobNnRPzvjYG2/K3aul42XMIKkx1vj2dnR5P3dYwHbOcQ5c
TDjg77aPXmQpL3DLgPuaEGpVBOVFvwlQyP+vEQiD3dtCQr0FSeE0GLNu/OYFvhrE
6CMH/0UiEn16VSBwW1pO8xrYGlI+CNk6KeGcJ1OYHWud/ydrwDnxXYqs8/WN3S/U
QNDRgLb+XnvhtyPvrmMVbuiHtSGH02xuJUGZ8xSt7mzfPDD2bcWs0VTpcRN+YZE4
1A2umczh3dgJzHywWW7aMhzKaDKB+MSKEVgXE4MFAbGrbEbrmMyN+sWgO48m30gD
73hwwmQKFxuyna2P5p8v9qIr3jHOyDYy2Ednh7RPesasy6feGh8zq89K8de9J3Bj
Rh1fcZkpXrEG/JuGQIixoCOOhD9azFWe6EFWHJfTHyDimrOuttiQu7VAn/nG14Im
IgNG2N72lh+3Pzy5Vix3T1OKbkDXrzcZC8jAIVpo6w8sC+jzO0bnlhC0fyYsSmpK
eoIWFXTmoZhDHtoW+7EIZllZU4Yq+QMxkSaRGCRO2Xbxv7tGWpDkxE0KhrRyPkCs
FZeoJooSp+LwddQALLKCM9emN4kRp9knICdBnacP7kTChwhAy0R5A2ldGT1mvf/E
CGFRNnyYCrTAjm7ft4vRCgHU/Am2EPh87djaNpRZrVwlqOU58M6bNQWi6O502CVS
21aa2oKK1u9bR4NrsCKVl7oMxRgCpDGbtwfimMfZ3rOeU/z7ivZvSwmxgCfjaZgU
dCqDopUgOeiZ6vOOhuirYUsywu51LVJvsNjteTtz/jF2K4ggn9JGkYMghvw2anae
dFUoWLOKfOvmcmaMKSjEK/LHp8lhd/xW0Vkr+DKoaCQmW1hsJqTSkEN69js4lP7x
hBJ2I+D+u4MMbozIE2qH8iILehlDuUi6pjTyI+NTrgS8zFD1TrEyMgKOj7O/mgse
BprHXfgt6yqwu95wpvcAbLXwei/q5R4JINmqf2uHjRSVhssBmMWu1DEMat+loBeF
la7OPG12HO74rRJPK3F7tr4cxtNgMvfwJLdM8RY+pIYO4e8/hhAqPrPuqxoG96d5
u1eYFlBG5STR0ibURuUtHxj56LKuT/jpi3VtnA3p2B7B5NZTov4Ur5WJtUzMzg7s
0NJbop/PuL4dz8SPLuZNIrYo0zuy9AusXDys0jnsM4Jyk+7BgRvZ5fJ86WbN608M
rq7SXBI0wm7ipktXDAh7m94RWghogeW6WbIA34+v6UqsHgJUQWVbAJ7NGc+pqyh1
3EubYaBOW61EWsI8t4mzyqaPXeXj7W2Yc9FnM7Yshe0T2No60zGX0CfS8kq3yll5
mjJsvBt/QoCTp8xO52aaZx4KnQrS54Pb+kPL1t9/Xr9RM5naH0CloNheLd3U5vZa
TBb2Fkd9+K0pEwtQTfnXMNB4kO1IQ9nc894RcZupq6FW+OGYRO6CtHEnnp/CtD69
o7vrw06kY1iK7Ec0Vbtw3ptPZiGuvk9Gf4iet4YPHhuPQRORKXJQ1OzdjcBPAwqx
2xmRnFJ7qOXeKEU3r7KHTmwRy/MgSyw/XKiCweDyODIYfKuRi/6RSki9znp740Qu
PT13gY5irFzEWad2MgW7EwQ3LNItAdVEd41Z1c1S6BcVJK0BZUzOKfTHNqufzyS+
kWwsympcL1sW+eDdFqq1HUMKR7lhLEOdIe2Ec4NfofA+G4VhisGJkZMso8nVCy5F
BGLk2SyNVCMJlWUVzlTT9MQVKg0fOOGKK3/mKSSUMTuN6mXDRwFwEuzIemxDk5Qw
96GHu9pK8iJqYTpWy/S+eeowZn3dh665XmVDHAp+hdmwvp/DhGYc3YeIWxKucMA4
z8VqD6p8XgNNQ0x9Q8gL01bRcxbvNZ4VpCUSQVr+fgwDc7IJgqMXRGmdUIj88J7S
4a4AIdArqs/ThEpm5kxTEPg4siqmqSGKiwGRuUQohUspKSdAm8AL+Evd2bM7ErT9
512+giwDu7oBnzLRxp97fXqghRFSuJMazFJlDEThoqHQ0UoTr4DJbhJawmUns+Un
rw6lS6fkFnhJA75zQbomRjlBIVhFvKiO6ZT+x+oeflKTS0zHM1Bbg8B+4NwFAyTO
STaSYdNfW/rMF6Sfl3+Xa+ROMRsv2VF8v2EoZXdffNyZbNKBxvKYvtN05/1u7Est
mVDYRAC+nKA7jqdz0hqjfNEPy0nd5sZ69l5W3RfbDwvRydhCZ3vfq/6PrrEi1Hd4
h3UsaAmbpuXWrrLo64ul9SXz846akbbdsTg1aDWLIsDcUoh09DIMpA4GVFt3zsU3
TLn6LR1qp29U+YsjEhQofYGtRJhUA+j6ijEWdONIAE04pcEa4njuzdjO6VNJFbIW
Ab4XD7vU6DYEdnJdiAR5sMoLQoWyMij/BUhi5twCJWD5jvPDacCNA8v1zhezoYLC
yPE6okta7TnZvDZqpSI7Dy6VBXiz4k4lAlq1QahezWYRuwcf5SYhvPiYXuwWdQJV
lcpnSuqqm9FwXSf8Q6iX5eWHJfjIw4/D3mqVkozhMKIxrcBMWH/17JoZBo4pFcIL
L9NSLnM80zdWd2Sm79lgxfp4cm425cQRbQUm0/XWPbC+qlNINS4gAO7t3vdjOyAZ
cfESO6qhvmhqrp5n7qxNIHTiMQfR1Udw/FuKiYyS1YbZjsSzJ/uZX47xXVkiVNgi
Dg/RrAnevzhTYLFfQMdYYQXKw6GCEcooaY8JSFSTF00yijy2PgRIl8K2XXwF3c63
vQZIme9Rye/E9ZS0Vf7lg3cEU9PClEPuAPvX9c8sthAjzJews+YM9v8k18u6gJES
dAxNCcDAjK+MBxOsS0K3ifVF6wX2IKKUjmz+cWtxmulxvjvoQz+nBieU2oFfHETr
JwTA2OfU8YD9WbRahCo2r5mz1TGVDR70Lx8EkwVar6OGmU7kT6yayzEWiZhpPrB9
Esms1kX/gOoV8ESZtTgYXuFCDlB4hm3Q8CtU+1GhJRT2TM8xBQOKwjDzW+IhCpx1
0kqyT8NzouLhtBSiSgPRMV5pnXT3+rxSXpj/OvNmjqLt4vVnMjFskNoIf8JwGwAp
v9B14llafEetjeNieCYQnjqI+oAblkDjONeeru9QUu1bNyUCJJyL5RAON62qgK2t
svpRIloLNcQs7aK64gPBfL+2A7xkFQ19IlecTr43ZkD6odtGSChPCgLTKdoRjg89
zhQUB0c+amkl8f97f8h1NZiqTTXDljpoFc5jZZnrwclM+4EUbF0dUmGBfJoDDNyI
rbM+PH56c4T3dMvWg6VNmEqUFVWr4tTDhglSzvOjobhzHCnpdPJ4x2TEgMbbChi4
orCleUfpKPW19OJmZ1HSWYiGDJgynhh/lpNVO3pLWawmtJn+xXusRUAjtchv2gAh
FSi63ZaoKPTtoBoCp1Laa8wLqj1MzrUwU0tYw1AlUuMjKrtdj6hIvSl5sU4uw+qK
SgKYPv0AHMR/o1zI2PZLyWkh22ZOaAibOtysngUaViwC1jEwGJuKFMyxUxqljkM2
JzP6ilE59VJGtkXGByekwWm5F7OfCUu1TpXSsYSK+MUW13ryaXlZ8mwLE+/LrE3N
h+q15oPtxgK+T/HRbkEfGnknNAjj66aZFE1arpX0N+Cw4Kh+2V4BkwQEJzWwYAYJ
K83zzq4SsbUBpekUZcuvsOHkHIqWDoDc7Jad8W0NJAe4gZ89bvd7baGd2lROC8VS
qUYiKaPiiJu7fzakJDMfniKCSgVFdyR7ef78zRQvZv78/2mrcttCyjfeCTojmGes
e872/yFZoTMZXH6jlkrxtGijAKB/3xcZFPwRx+1G+g3nCxRno/ddjgk1IK0SAWqJ
+T/d8luxyZ5zOegwq+aKwTmb+xvIJyHV8cv0npCrwpgQ8Qng1h0j5Ml2/PexygtJ
9+n1y5iKtnyLRYXQWX3y7T06e+M+qInYXx++i0imxTjHE9xyv9jJMBLbWBJM3IhY
zxc3c7IHTadtRzoMJWncZQhnQD+Hx8AoyfC0OJQ0aPevMbK4sjr2vPIWEFtKXZ4X
H1JDOt0ms95997907+O2kAW6R+IOkkdl1mZCnC88FULIu6F7P2mnFYMxrBf720Bn
4UHEjcwjrslQilkb7b9B571PfXFDn7WcTZYM8JgmRNfl6QSzobz3XVbxTU2Dy1mk
0GKhW/mOotID41SsaTF3YgTki4NNWoG8Fc5Bg5YyIHmfktbbFXwdyrF8jN0JYoSr
VbHI6cpFod7BO+B4hJsQy/L2fn8ps3nyTS+HA4T9zyIWmGcxXgMgIFJlNeii8/gy
uRsTLgEr035bjCw75XOBq9wk1l0o7dNAyr8aVn5bS7lHwXcrY6iBwkihH+YVzoL5
WY7oLEB9Z6YmxFv/shO80k8evrNJCm92/OTj1N19nKKcYCErUgvqUmQgLD2NT/2x
qcRv/IM9KDMllpd7i+4/P5WSW2PatVW//5p/W9+9tbkb5VlmWH0N4TkJnb/8xIPO
ohNlXsAj4j25aIeNRkpibMo+y7fSZLL5au91O2aHJU7tehIVSYRWQR9kprt0ZVS/
ZbbM63NDHhUzlmijjBK8GK36HBandYAnFJXIDrAIZWITgKYdgFeUuWnhNUzUHIjr
WmRldRg1R050gIhkmTIL8OuDzv33gBfUDLHbUfLfXwBsIRimZiuQuUeUFwz/a2Z/
XXd38VrOtZacKqbzrg6OAD47Ert7KhpBhsCFdPEmMOx52MJUUIINlnH+BEYZzqfb
mcYifNi1+ig5LmTXNG5jVsRqGjWF+Ld1RnPA16EBuk+KUzlAQAEPoe0kmBChOnJF
KUzbb9A45YQ+uNGQY2lI9ph5SEsUBQq+UKB0DW43WS+L4M37vpn3MHBHLVLwF0IU
VwqI6NJbaLEvgUUG/9ZF7k4DqYksAe5kdU802c4EzKKK/oZnZ3TFsGhbVv8Nfdzx
rFi7D/fkoUyLfqIGnT2e0lNYb9Bt4KpEeLaGBKwaHN27EYJtU5wU1kThmvOTpDUT
3VF31oFHO9XXSYnl0hW/OPab5LVtLog3Kwj3CCMEohZbsoO/L+PjGulzqAc2PQdi
BcgXu040OJy5gKWTIsA8VTW3gSdW4NpxKyOvFVAWgRHj4opqn5OfBPOP4KMbW99J
qeu54Trd5smPbNgiaOmeo3cdVUSynJlQSPaaI2loB1wxnNay8UZjY/DdV5UtDJks
mvi6ijc4PA1aN9qrR10LcsQ4/N++v8xMrPiqmJS6qX3mvCV7UQDSYs37CH3B3oop
asIiAAdPaLjU2F+C+jxo6qMd7BNpwuxiyfMav3GUra9MxdLtDynx6rcL9DEtbhxV
/cB/1ndCXI6Mxuokv0FPvIue2NqbTmvVhHBhhv+PeqrXJdq2fg5al9Q+YYKzX2x1
3auwsxMwmF74OoK57AQ8bPcnQykNPTKSawxfSYwEjAPDZTsZJJWYY2I2A+xlOfrQ
j2w+wFHnma/mzTbwEwZO4DTyHtR+hook8GpipeMjBHsats8yVh8dxR6kfKhJ5pKy
+/bGgK7kqLdBVHLs9uymKMKrOuIWqw2SVvgSjsrqLPSaytP2TP985Pa4ypvcj7E/
0YklkcZ+GOMpxFDzps4SMTP7047qnyWToJ0kPy6fk4+aeqMfLaGdiKziVDRsxIAh
8TNSjBe88V8VOqCxrYygpB2gzMXBOSBqcCtI34evk78gzUTxqkumFm+iPWMHMQO7
kq2u1sRBlWPPbQ2b3Se7ACUYFibC94aAO7fDvaEClRWZRovSMuqFapTnS6V4DriR
telZBP2sbDwaW5tK6Lp9o09eRpAXpECC7Fj6Tj4pUepW87iNnthWqt6cOd/EkCLr
LjYscYrg0lhIwZvLUYwNz2bouADxhi7gFfifTogHGb9ujpR9xE7wWIzhANKAust5
Ooc1tQEWtSR/sIzsF6KfMcD9BU2RMe9nIhpV+g2WjU8lsjEyc/7u3rALUf4SdP1S
iX8I40haJ96XE7/v+Ry3L6EByql20QExL4RiOdNDzXWXj6fzzBD6XqsrW7SfkK8m
paEE24Y55XdCOBkAg3NnNiahVpDwH/jztDpkrRHJW9MHPnEazdP+5QI+p1JkR/BT
fNR+8j8mZXJE6vTIz0qq/3+nhRMWz4sl/I7jmCJ+cPqm4tjmTovuT5TPBTflZtci
+1I7cMrJSx9BxllgR4qghDWiM5QBu/6tssOxNitrykpFnTKqNBwRPknISp26Zn3R
1nut3MxRZVW0v8mKAzydnuQpyT6V7JNOzr8uFfxTfc0bQyv+B4lDlQyu/91y6ajP
wCIiV1CvgtgXJm0WURsmDfuZTGgKANpir8kzmmND8LD0vHRJsYgZbR5v1Z34W0Ky
umZo/B9+5ZrW6IluSBTrDLcpgtBuBmNr70WBfBGovtj3n5JjDQ1n8uS90AdC6PX9
qQSIQRmXLAdjAzYXmFjaK9nlzUZtA3YZsV0flriHLSWFptMcTZgztnj5rEajJx7m
lfeS2QLUVlhnFr1fAIkhgOw8T6aP7tMvfaS2D6zTT5huObQ7XIlUxQ37HTeFfcNU
ZWcmp9/0ZRaaRCnlUJnBzDiHnNqUTuKFC4/holC3sVxcxY9rMp8+H1ACDxIHjFy0
Jdrlla2yPBidqWz4FEBBwX24L0TFhyNBrBpVcOQoXQpxOe0fepSAiIdHVJbq/Iym
JnrXJqnO2Dzh5P5SkAKrpRtvvFcUnISwuLQ6qt6VBALvoCt5X1rMrTzvGFodMG8N
otWTsS/h/gaDRI+VbF1/u2pD8/7YjEGja8wOetT04U63oeeQazHsT9VZNQl0b6Ik
wAlQD60557CQWnPwWBvTj+EAKjiDLHIG3OZYqjfr855S02bJoonb9cRhUY9arPEX
H13lttwF9i5zm3KQ4qwJtd4j+URo2oc8psGu/EI0xVG0SXU75ZSK2Gb4qukErQ/I
Nq52Tm9hDi644uhURuVbn+36UoPFB56TTfkiuonGPxMMzNTw/ilWno6tKiHIc8ml
AzDqalfAVi6mY8Sp7xn3/8yPnEtwsGHMCGQCJusa5TuYPghqR0QNQMHrpbe+N0pA
Ewr0zA+w7EACCom6ATIV37/Uogs9z8CbcxNvBSYX+1lExeblvIIseeTO7q+106JF
H6EV8ExZgu8jRvEY8zR6aZryIA1tkjm76x71gyaZn9M+weS/riB8DYNwTbcD8UzX
1BqbEUlR7/3lvzWvgT2lxIVQ8HZWhpo+lbUDcpNu+oth7q9mNfhcgU6QLCusYXbM
nlDE03hu9zA3RH4R/3pQgkBQbRLv9KiuPYZN6bP9H1g5rjqepxRQOvax7pcgpqja
0ul+x7BpCGbjldqrYDpUB1jFcmYxTydZPmY64aBpeSVvDGXbgP6CRNgk/LqPSF9y
80y5FioCKPPZHbTh5eborl7CTdDX9Kr8cP0NNc5aTaKZ01ofyrgrn/aXouGgrIJP
9fH37bnc11NMW8kUzsxtfgvQJ2uVAxGFUZ5gr0RVeAM/C7xmbn/5Uno+x9J3UYVB
ZZKn8FpG3/DK3SZaluv5f0DTUYCKfSTIjvQF3uIeArlUY2pLV+wz8MSUurvGh/h4
Bt0Cdo+AhBwSgPgL7PyiFCgxitAeCl1ZGUkegUuDWTOJ13mQjoxIPICpclXjN22d
WX0OhVUDBH56aV+vDVEEQ2qJ5XDSYeawhRBroKsxebN/vC6b3pRq5sWF8GWkP3zi
ev/1oOp304WPSEDPZOI+1nS4c6Cf2ngWVonT3DnbMVC90Q8cl2Tvrg1d5ZU+CKF9
nDaorM568RZuK6b+6751hsUE1isGvPD7bRB+5QVALpK7/IQmcVt3F2pMYc3IoY1x
/vYdIbrfq801vFvx7odOF7cka9PjFC0D57pBN53B0oKjcqQA7NDpdguSfmJCIee4
5/Ly8A+g6LlQsDYqt3IGkPRKibBIqfFpH+niC+mhYpQAklXSQ5PxjQ2Cy99vuXn/
p1PfYQXl7BkcKFg3TR3DIa58F5covgV/rVedm7bjtIOHZupqrfMI6Q7P13dHx444
hqTqE0skLKgqHLMydsC18LZA2Nf4SFjMLS7raUocQNJDhLIvBJxtfMhksszNIq4r
CukK5HoPhNPs0Ri4zIuNeLK1sLGXUeZdUgJ3MwpL/IxoBy+SK1qzCKRESeX55dtF
pTrXw5n2Ch+OwCoe7UFrBsnu11pKKZtwMYp/D2MaWFVnTg1oMw3fovYjYILCl+hG
EHkCc9wARm6W23Zi6pab9oD0RFp9dWmhoRwlN7NqFXs9QHtxM9mJkjtrn/ZU2G+g
gvkxzgqrmSNc7ql09LxTzfsPdowkVPVu0+flc89EJxa7Z3m6/xQsk8Gq3gUzDDmj
As0h4Tleu7XYzxjj7+E5dwCZnBNwZy5neZuPatmeAQUmTXrbXzpZRhHuRI/ePAD4
XT6U/YiCsfj62ooqtwZHX9NSAdhvpBXQsrbicKRcFmHwrAv0ncdwXy6jpgVuvLaB
GUZijQkZ1U6yj7sFr0aJp0u2oBXRa/zlqsdfzCzaUMnMwkbZC0xzTJwyRQaNA/Qe
ajdtOOnVRW/hZg35jO18p9EMqv2iosQSIQ1VD8TdneJomoori8zJj2gmuhcRCHNs
9GX7SJkK6odnHVN5iieCDCuMCqQ/mn3ferjXzWkulNxPCpE4mPStM/UHTyzFJass
P+Kz/H19s4djh1MGXTszYIwGdQfx0BzKhvwXzyU/45bRE22bqJsw9sM6TRwWzZ9Y
pL24+meE50eXlECy79nWQlQPtBEFQqe7z1qtO+o7JnVPwxhMeDPaRJ6xC2EUme6T
zkhk641h4CjVGEoIznwjVsvR3ZBQYXD9PmcnDdtAz5gxt1hn4IMugAWaUGGG6A3T
v+zGXHq9gMpyPjDwCLHhkFsuTmd/qKWhiHQJ1tcvli9eo35tyInZZfyW4zMQ0I0w
jepiBNpwgQ0Mi0fitDrPPmZ0qwUjiUZkUJulxC2x3BneE13SQd+IrNZQv04rZoOn
51zPvoOiRFtE/o8hdN83hNtJjn1w0YBNx7OZpuYc445LstrvMR+wU/ADENKuxsVe
xCNrMpbtQ5wpJ8EtOe9zGMToVqGGSyco6jRd02OUxTZNeRC8aCLrV3oFm5jmfATL
JhMPI+ytRvBk1aTNK8Dj1jmUy9eNt3G12yuMSO3fkQ8CCcuIjFaz+bZNMDjOAzje
yiSHQmhCQ4GRl3O5/Jxp2pK/jZrBfUOhjLbtmQm+NYJs9orBlXJbE2iIJxut069X
PgJeELLbS0MWQs6M9Y/ceon8k0f4csbkpyRaEj2NGKqQlwzc8bP2SgHsO6ZmvaRX
Ji/3guyVgoFLaRSDJJIWmdshg4NIELw2j/hb5x4IrtgT0J8ZQpcEFYNcI28PVNIA
skgfjBQEWwaSvDUYXdso432+KbYOkrd74Z4XnWz853X9zofXYeLj/yP3LaZ+USsI
eIJMVmA6yHEy3MKyIxj+9/RzRZqM4mg5gNEvN+IXEFq/rRPwRvVrZLbMYHz3kIY2
r44sJSih5NayuN0j42OF9bnVSnMXpxto3X2TCGn/5PA4oq1Wl+lwj+G29YWNZYL2
Va2lX5BC8oRG0HYnZgzKRD7g2YaATNrOwYDjhAY9T7+fnyP6o2c5Q6BbGy5YnM+f
wK/hd5x9q1cYsy4/DWCkYoJ85mEJfiCYyPK+UPXNjTZ+Tai8LfOfUSlihzVGDs4V
bTyzhKeiaWb+ukme921vhVTlLssl7Z+ekh17pttJLJq7QKXigiebWip36wkzCCI2
3jS4FSTuQyX4JD78EJ3m5uV0HNT81RU3pJvsOSNnyPaEdqZ/7dCRC6Gc6xUzzrOV
rhJpBMQ9+uezIDL35K1D016ACTMhplA7LlYi64o/9QQrsWhSKcjbt8mqRcTzdSl8
cl7cy3ExLzR5vvjZ+hiPJDfWian0uCulwXuyonCRkdmBMeNxsf0m7q/oO1pTxBlW
KyugQFer+eK9s4/sruqdzuoY7GpAORQ5hHLNshN+JRcRchSwYrS20x7nAxnpQnEi
Q82DfqczbwISwlST6LzesKIm9xFX88QTA3sxN0hnW9twASvr4iLhtnKvQ/ROaVoP
6qJaI6QQOfMliHGTzEGh/T+NP9g8JgKcfb10Z/N6RhFWzYF7VaKT1EYeQLQhivzO
wNkaBAxboLvL75NC5HdDoTLbgcxbljGDmY2f1cvDhCSgRRg1+sGkPCCkh1gH8P/P
z6wDdcWIlewZJHYd4nKtvARlhLQatZdDQWHy0RMqdXHJ68HexaPhjlOx5SH+JDFx
icQ6K4H8ZmYOwzjwWVBF/7AyYqilLsbtiHDVTjSrHELemfzWK9lUOuS0v64sBlG0
DrOeeVmcz0BuQ46bFoIgXdFkX8OOcLPy7ndhyelg69Wi3rePp033DncexNhPRM/R
EexZqk7yc01gBW4WdDZ/UY8Yvfe1XVePYTREGamcuQQn57hsY7RngQjTofnRAE8C
bl4wY+NaVb7klIFHFKBU/8klE8nqXzPbsb23Y7JbUvW8KYYa4PWuVM0irTxxqoH4
wpD6+vCnh+6uxObzIHRoROBH15+d/gSoS3BSl35AM5CvPt59NBLUa7o1vCNETv8i
NzjxQTyy3aFHwkSOTLc3JPN3JbHKbM9muySytCmPX3qJR0DDJ1QZNTt7GehkGosS
nfyjWIM7nDEBYLkcYhoV1YBzlq4Zp/SW32huIv+O8/cDEBdR8rtRFFHYS0DPNLzv
MJ7JkiA6ZeTQHVeRvEHHvv+E6UI4Gz8E+UwovmxUgi24NeNfKaecse0vlyDbwnrZ
p13+FQwEZ45brSNvM9RHX+yVBazc8dMUmLFQ8nR/wzaI55sbL1UfmLHftwONrBsb
qScoMQqnXuz81rPUSilQaSeAGLigg4ZyY3jepA8lhNEDZ+LrRXVwNO97pPapM5vM
gNf+tdrEryZjD5KESKD5JYy9MiUlAiJRf6CKuiG/dtFlTw/LwSEic/TOlCWtC1/2
I95gGuGZ1jUCw80il9DL2e67jhgS9cInGa0Xh3wzJv013SsSrQIVjn46xxs7GKK+
PLS45uYyJwFc/Up7O+oswzJ4LDIGcbsjQjOdUM4aL7rbNHJWk75qn08hqQMV3I3y
/WL00Zbi5RaQ47k6z7TXiRcsWoO5bGNayXbH6Eqt7K8YXA8/fWCCYcJcksSgG7/O
aNNHoNnFJn7Qkid5SkHSzr2li7/SlFMc1wxnNWXYP8Mn2TvtQuJH8Mm4oyrx4Pk5
usEu6BNjGgIHj49DxyCItV8mbGZjUrw3+oupVcYOO8e6/Bxg7fU8viUTPf2mq39Q
rWrCAq6bSylwtu2YsO79GW6v65w/zRlkWMfZXDBTvSVYLKAmfkA3UCIbhZ1k1EpP
IOEcotToq7g014S1drN2l7R6DlKtW32u2y3HuD9pYpktviryfqoP3eIoNuJJ34UP
P0/CWaggVug+OdZhQ+o88rImO8pFK/Gwz86La//Wdol0OXhyp8qAzzQunxprCunz
kZXd+ohKLsv4UurxnHitTTKNSqNA0YkQMQWF6nTmfIpKY/r3a86aijwEyxRkwu9P
+fWT+wy+vB6C6kPleyGdDm5j7Co1IuRML87sIWmzYTObzdQ6uFfzEJbPiTdp79jb
ECMszomtqV5auZ41T2wz51UGCgXSxV9F67umMSuPSbCHsPvUVtYlmUTDr5sIDFmc
D4qjY+NOlwY3aPrII+KkKRvHX8pFEjT9kMePwHnzMQKMPoOIizcCTylR/1jYL2Dp
ADS+oeqA12yXoxv7jN/ftk0FqtuzKUI6rBlSCtOZwfOOrL61jGLYs2KqhRfrc06P
NxuiE0VbE/QpfddAZcj4+kv5EElaTKV1pnIEzfp6bpwabmJY1yKlGS4Qtpgz+OeV
YeGF8t6cDa49l41Cv/nxDwfG5+F+zMokUSt20Edr7VW5m5zry1WWEdvp/gXrZV9u
HIEZ2Z0yayDrhMcM/2YKMx8PHHj9/nPEXD7evIml88oWrPfg8QY6CEaImr+GzEE9
fc+ve61RTAQHuHpTVOJherZI65m+yew0yRT3/tWln3f19+D6jOttOCmaI1VFlwB4
PLFKYJjUgZ84X6atiZEYAFM462SPaIi59JYsscpAwHdk162krg2ttEdXkhQNjZal
V27q6rJPcPmC+JBi28CK+RmAKBBscn4v5J9qQ4L833QdxOozH7rGrDPv3ZZNvFK6
yv9KELkm0AMXFdAvbchGI8+aEp4G5wGC7cvTx4ElreysOU5iS1DlYnavqKVxrj4N
Bc9mrEA5S2tsSQz+lpG+CYjJ6/cE7CWYnrIyv8OfR+cJJXvFDXxWG+jEzYdWtkFf
hDVqUfWLv/50Jj5Cg0edzrriei+ZOFnJrDU6W/Nitw57nsQXsfV+N3K0uXVeipzD
0ZZFE1WjG6hets8vKauwXozIowcOs05CfZ5LkJ08+J9efeqVqY+oQ7QuwMhsx2pz
lhYAu599ZFeXDF+7kUzXDLfkROBA6bydkFHTpCAUR/HYEGTx6G/aW8aVSiyfS0f5
GZvJ/2H9Y+xI2+sLZYMjMnjyn5/i59/acSeM2sUVkqy6vb+epCTS9OSt086TlU4e
tYWUoZW0WDbHdnnKuBYhSCCK6wSxZXXF4REEbi7c7fGxFNxaNHK69T8GZPnrS5i1
BNnAzstZq1RFuh7wCgTkI1VfO/f7DzdN/rAO57/6vfHxp2DcedIVWYVcQKELeDrX
+O7X/1YlseH4exqxZyWc6bkFybmucZnz4tV8YakFLbsFD5uFj8/FihigDWwpU8CS
lDUBKbY9MYJsLXcG82bp8SUpjPCYBOPmV3fFh0eFwBN1FLyOtJFdwyY5HC4FmVH9
oOJYec4WI4ga15QvmY30DMJYj2Onv8t9PgzVMVWLqu+TCu94IKodFZFvvGxht7iu
21CJRZOLlV8U0Zt+5uuiAmOrpbfXQ1MHfFTe3DAPLzRRpT52X7TEBSJmvyu540lv
rC3VBKAqpW23QpEz1LAuEolDUSMsZNh4hpzMXH+aUBBQPZMlMKRWd4y/N0HzOSYg
lfWak3dJwhlsgO4bNAnp+uwHvaKAZWd9IUxtwGhyukRTzuzRrPsBC3d8xQqZYkqr
xB5RQ8uGvCpqzo+tSqOztclJhOpQN4OeOIWxvP90mfApvW5n+CujsKPhhKtVlpDd
r+kGfy83N0czzRmMKhYx3XFLg8LRfJCej9jld8vkJcYQsS9eWT3+1INGT1PxW/8w
AwutIzMvmqUqBmBeKCx6JXp52f6ORUCv6LULorVOYnQNf5Rvf+ao2T1pZDkPjz2M
H4eNONG4K6ZK2/f1hCcTgllvv1WIIo6Ezzti21+Oo3AEJ9lB3uDtRTkyDzn6PMw7
vA+v5qcn6n69EOFWNYg8Q9h95LVoT73iqFKbhnSta5pSHxuakk8Wg2FEvXxYRkgB
r+cU3ug6YR5BqX/mwfVrJvscX0PZSy1xIpdO724rRIb4ByURuj3uxrftt7uhHPgH
TbGA9df6SilNDsCE4lBKCz/Vlru+BtyGRCaNGgRPBjVuQc/NVQLHOPPGsqBNZFXr
alVwEG3zxazMhsqNO1/1YlRFW3b2SP4X/ouephUk9rhG/1kOkpQ3wJ6zWQCvlJj5
L+3W54+jN86UO5ivGwF8FLsQ9Dya0jJs4G7KT7yX64vjK4YDtlu4dJLuNb55Ztdt
OzawsuNNODe3p3wsmGfdTzXHQ/78bjpTism9pERBd2l62q/gV5gdIPdUIkXyHYRa
5y5vjaz8h2icz4PS8Qw8dYoxFJQPO14N8Pa5UR0NnBwG2FeTunrRiz4oWc62+4o8
3B1Ymep7zUUQ22dKNTZO/FxJlMh004Qowah0oJCNmaaou1LJW3ox85vdQM33tsfQ
NG8tltisnZXgwPycA4x3qaFCTEm0Ie6o7UMKTWjxI34Hk9qI53Ap1Kmdl9AfyxOL
UoGknOkZtM0gzRGPGR3+v9C0GzIfcZxbq9QNdCvhlW802pYtrqo9Kds0+OYdk4oi
AErH9f5EofgLd+6UCpagbW/e2jJao+SoFTQ5kh7NO6QlnWfXAC/EyP7NLRqk6ET+
LEz24IFUibw9O8cbFpBwojlgA5VuNScVKoSF8MLZEMgrrb+HoTb/zJ3e9T5tCzQn
HZB6EZYafqBk8gbFoxd/Ig7t89QodiP3WG0pYQX5ipQYA1xrHG2DceacRQoXjEOG
oBxRd6yuMD0/Yy6t2Cn6Ym4FlYi6/fMrwKDQ5CxoN2xGLSpvFyoyVuANNYO+uu8R
W87veu6J6IS2SFgOa7FzZ0CerD/WWX1nrGqQmQr2oMVYKXWxysZdm4ali8wgQTA5
6qzzRjXjcXTrxj+HCu8L8J91DK8LtkMSHsU9R7YsI5x+7C79QU/WuPj9M8NVoO2v
/gfJVSBQka9J9vHkYU1zFfBsWYDPnWMD8ckBq53v+pGBRJiHYFcuvS7IxapjbyKh
T2UlBRHIPXoErnONt3uZqfogVte1NIAsKCixNfZgV/42MG4o561OJw5+JcDsyhRg
6yS55sO+DxNibtuKJDLKojPSv0tJRO250QPHXpmjGhaBI4V76png02e+9f9lJ2h0
8Isjsvp715fdAD1sKT6DqMUQ6Jl1Y5O4c66Y5bhmzjdCg2EIfk0LQpuPWUw0MugO
r5esZHEJ7OmJUYX+prTcB4kxaM3nrA7EpU/hr1LmEjI0Qa2x8Dp6Ed/O5ZFmAo3a
v9fKupZm23k9FIL1It2q7biNJ70Y3aSyPRqP8EvurKsPp3y3fGBVc+bSe3jv7iR4
Uoo49pm3VxSuipQsf/mWvifeLPJQR3C3o3cUYAG400Pn70oS0V/qjlAguCi/Ygqi
f9keyf2HrLuAUnoYiOBE1lQDX1v+mHO94LNIQPw5xezf5uFWyGZufkhzzeYKXpDS
0VlO+arBV9sF/kmeBSOg0ldYhHwVl0/ol+R2EsSdoJhTS/u64ZYg35UmLhfF4eTs
IwsUL90y9238vpP2OhdxfegMFTW+D273DTXhn+weoW7dhRoINDVNpuH1bhcUtKHN
s2fTiykIYxIsAtDokEQbmeNeTKrfVc52G5EanE9MzGFL47oCQ83E8bW2PcUdLwEr
Wkc7nfxct9kVESz8EP8Bay7bR+uqkVcvyQmVRp5Kuzm0n5l2RlMHGhF7HIo8UEZu
VVnXpOYcaEupt2pWttaMk6dtSrpNYPfZO3yFgzTS0J0vqIHPCVCGx29ABkMUZlKZ
SHIB/B65owR2bFXX4fxVQEwfkC2WeGrjJ7aBh7agGnuxHuWPPYwAXd40K3BBESi1
s0y2Ux6ExmRLIlOuPSmVRKjlXcyTIWYJI+HPtmFd1hIdLzssFKEFbwUvvkTp4P86
fcPVNlsvdKHOvr/8L5cL5ASYiib1NSpBWviwai01VZr/O7vCwk0rPh0Y3Vt4EsJ7
kSrdenvvtKsXLNNaAEUeJNo0LQHr+L4MKiizpcVIqYV/PrrD4SaWq/MLyEMVfjBD
yfaYCXZM03Xk8GiJnE7Cp4p0g38q/ynRAbnlzCD3+WsUakdAK4pwRvQnptHkCYZ0
n0I/LhZk33YwCAfo+w5RXuUBEQm6ZAkIfE8EW6EZbX3VV0pg872lJ3uqoE57IXCV
JqwtkJ2hhjx91zlYX/vQUu11LukU4RsH8ojKsL0G9FxsHIxDjLK32wWoUxTWVrfa
sI4gcGLyqcNnugb4eyyLX638e+8ktA1wCdDo04Ksrag6xAHc993rP5dZCxK17JAx
2VhLtbgu98x6NaoUcfR6aQGp6bHJ46yXQo410XM/pFOfh9XY+5nkbMP5FakUWs/Y
oTCy3Pl6it4dJyr37Jh2aFX1F/h1N4ij7KZvEgorBPrgxEto/WgiYhE4DpeLTeYz
pBYf2C6YICBN1aj6RR8g9sMDTF0Q0p5gqVHrp6xOo+Jc1sTTqxgOPDfv9HLjlIZi
j0w8bYCrzISV3dscUTPsEYW2tvvBoibtPQEI8T8A5RjY6buiHOpRG2u0DEs8cg3Y
pOyBCKIsnhiz5psI3IyfBuTRuOilYG78GZU/VQDt3jqkdlAFev0LNNYQtA6JTq76
GUPjmwXlcapMMr9Jz6V6GYm56aY0a9SSV7yG5QvLRyeqEDvDUp33c9HXwsgfO9HG
PRxN8kNz/l3JJ+fnxiYA42bfyur8LLdFEpyO3WfO2dBZweGByqFWWpq0YoS8h4q5
mRLju+oydtiaDIcwjugZUGEsIYbV04+rBf6cXw2rrD6KQJpoAXeoI9yZOXnLcrPV
xiVn4NCAP4LVIHTY/AU2ZRi3smUcgzy7OuIbUY/Kq3owVBrtLXEXGo/5PueCTtL9
XVlht6ZrCORLKNk0jtivRMRpD9OiMyRgowIOYg4GmqQWt/M3MHWT2b9U1Ijvqu71
FMchzlfvDn9lAQIcBn5VVEN1lPfoc3HBj8Am3zcVq0SrC1qdP0WxiyrsmnaYTiH/
tzxvqCoD3mwSIq1hnp7k9Lwu4mC57/1s895Swu4A0hn2E9V6EKzXD194xE/huLEH
cR5GTCyxf0Mdtlee1p0aoh7vvPZ1ho5wl5epspvimWIygu2WmogCoKTVXEJU+ZtR
hYSonNQPb3HHTf/DyH8Y074DmY+zDDp559jDuGIg5yzWZGMYmaQBw3MJScVH56+j
wOZS1omfTGcObiJACs4uucwkK+1j1JlBLbui/aSssrJ7sCrHEpaDF+Drec93XOFJ
sFzseIIznQ5Y96pn8Vi5e7tYZQuHb5MlJuFem396fSRsRfqOIUSBUC5kVrAd4l/0
3Xu7V5qgDjjTGVrP07UAlgEtbzIvdo2a7AD6nHDyGOlyiKoPbVV9OkDGLTw8N0D4
I6KIkwmUmkYwFTzYXVKHE/UW0YeHePieejnG3R+gE/8jECyq8m7ywesMtKl/d/8q
1jMMi3CximwKpmaGTeWxG2E1p8PuvhGv0H0i58QHYK4HYQSbNCLcgcGZ2liQcbgJ
tLwXuNuPujtw8kF8G3M/qYIFxn38hgwYd3om+K5qLjWMQ0ZSow7SAUmsWxU1k5yR
6Xj/Arj/dbDC4vPAZzwMhhqRYgaV+dkevtIN/nBRztJ79iiLjD7S4pwPovnQXlt+
r/2C1iqxTdpqeIkWhhUmbVG44TTUxwKMMvNJ5qWx/umbV7HcP0qllTzBmC2WCpCI
Q3l6Ui1g/VV5XH+xtOZ1YHHMB3VQMkTE8/x+DCfWEElywWUDJw6vhN0pa+HacKXg
4QMI+xqAQoaU6pgFSXYqvHaUeC18YdD9W5ugjeuGOZksEXTF2riXb0SVGpm5+LB8
CYKRIlnFNOdoq4L8WXlRalIE3JzKFGGrlfL9hkr12yMVGQmDyV26JcIBkvYJkgRF
Cr04asPJn2D1mBthVYDdfZ0W8IsnuhqDMPzBj1KnaA8sT4tAzE3T6tNWe/uLQoGm
kLf88hfeVcn6mlrEdl5BDcEI6kAlbLItg7CHXTE38OagR2H37vxx/g9KRdMzHA00
2VNhjzI78Mb+5kH2FegIGN4T+VYoOR6EcW0b8//9olelEMSoBYrk+uqCRyNPjKoI
Va4gcYTRwn7pr177teFvW8OpfLoGneQmiSerNbuKAU4r0IqrRGFEWtwc0wWt+1hy
7Sl8Vh1a7U+xDbIa7Jz9cjKF3nW548SQGcNypBc0jf3wsc07Kib5jDA3ERfaD2sF
sNVXHhT+GwXp3iVVI0wY/bsyUsoHeym9IsJ1mwXbQQeunmqJ6M5cwRP7dUg1+HAT
77ZDkgd1GG61lumRLPxHexB01lvIP8NsKVUpC02vX6HznJYBdyveyGMmDbkNhCG8
3IN2H91oSxaQKj2B6FAyzTJaijcG35vl6vdrS3/nJxfgoPTvltd/e0AmAMRC4Ni6
X40bVPdYAEXu614W/pR4l21P4ekT38SPKG4l9QFvPRZ3yytaK8RKvrYBkIhCFacw
BkQTRY6pGm2w3mjIYP4v+eXpfemUN93PutQ/pTMfamkVkoojQW4NMuqPAAFu6aYN
BKLPY1YF23NpXhheNZyGewGXP8p3kbJtYvaAc73Y5oMDixatViIcTkVnIOJlZx0o
wMHreSgT7zQlT5HqO8X1o3HpOfTYV1ZOgGBVQeNvFWxuGBA3zwjWTU87Cj1awj0f
wEZLc/ohtZ9gZPnKevxw55dwkbEzH1/qqI5nAyPXhipkzE+59H/9DVx44NLM6XOZ
rbAiIoy+9lcRkJ0Pp692+ioDBCN6q9y5TupfL3W0zpAml0NcK6hqupZrSTEhmSkT
ox2l3Eo70tufBwF2B2msi023DkN4Jik/nVia0q6yylQguwotgXvFBR9QiwYVr3oB
J82BDiP+FLctXHgpxKMDA0ZSaTkcRNZlmVTXlWor10Zzacgno6jfH+2xUf8L4M1l
fUD8+ZmUDr+jdPDj79ax4ErlRrA3dLhvJCj8PKOhUrebsltvAdU0Nm11wi9scUiV
Ib64bNgcxhYKNFGteqrJa7r8ZC59+G8VbJ5xufUDokWz10IDoaXdCu8k6MjePRm+
S2M7cU25Y0IP7duvreSeuEyyP2HX4yfLfw8RFqUDaJPWY93com8BiPD5bFf76vJ/
wAdUrYnZgovcSGGXV39FRIBqA07LvTzBX9S9R+/aGbcrfiZe2AnDviw7fzLlhetq
I8Fxd/73pyzaZev2xpf3NPYsi0Z26Q11YF9dztLyzTVzrJwDeCBeixxGyoErmaVo
LtJz202eEXTdATS3wuXcvfgYK7MqcFeaK3YLPPrwo8C3V0Rq1DmlpbbsFtYW+fQO
1R9m3Ig/8Xhf1CbQH3YXMYTnaFlz25Lt9nsO6G3OoDl3TqxS/9kD0ADUym1fU8XB
9DIdpZEVS5W/SLdd+t5jyX1fzrsMm6sehBUPjnbKAcu2TFLJ5UWCVN3SW/Lwd218
y4T2OiUop9RbLz73g9MBIeR2/8+aJxbpEfB/Zkj549YwXzsNl5xEI4xGhpCU647R
ns2KpVAnMdVuzDAdfpGwoRTm6RJBvSMuVqe/IcrX36hY//crOC3bfhNm6YzqHs3x
gyziDmA3h45SUJeMQNWwKwtgG3axJpmZkjNrAV+yOzD5BqtLKvvFFJIEyfcILYuH
ZanFjzwW8YhrGvV5edHboWzpvDeUlubXU9Bg22QpEXV58UCCPY1vSiRzqBnN+k6x
9ljG+kGXst0ndZ2vr7fUixrokcJTVRDGkyIS+rWyTOMEE9xzSffAAIjuPbUSrQmh
snJBFVtLEWsoATMyuPYJWO0bW5su8+dHpnDsVpHIvex0GU5687EqLgxbjGehL18o
qDAX31YamDNUk84rSfMVvZKSfES4iY1FDE4OPvIoRalp8Pql2MKauWDZ/4c8UAt4
9GAB77WJHRwD/YxxWxOHVHkExadH1klcXY8vD1XAj0TPRGUjYR2pWwLS+QwS3mSe
P3ldMZEhLmbHDXa1LI2cQpqK/M5JaoQKk5JxlQR0xX11ouOhL+5uTk3EYxvYUx+g
UgjAvWvyB0j2v11OkILW5HNE0MUhGutOtZ7FEBQLjV4aq2X1iSf4zVTLYBN+Bsia
SZ27+uATjyQNZ4/CtzV76eI1Fdj/Wf5kT5+2qVdo+bxNF6G4UCcnT7mAnX8uIg3Z
utcmf8OS0dkPvI6z1vBod2CyVu1qIOc1oQe8nbPGh1F+YEMbgi7a3lrvAbgmIFF8
yvT1flQiogQpGCMMVM6idvrAP+yYZ2wLIdl/HEMmXUaIm68Q9DL91TaI1T4BRYNy
A8q39VUyMaSPcreLoSk8GxVqiZ5Dq8M/F954yPINsrE35En/1tR3Jgu+A41RghZq
ZObpwsD1oh42MgpjfePw1xvSl/Xs6tajOGXC2/v0CyokHXkWtfpSQNS5qrZsyjhQ
Es4KG5LsWMLHjunB4gZMorQzFOQu1OJG4SWUZvGx7bODzjZH5gnPTEqOYnvy6z3K
fMpMAhHElwfKqwJrRoxQXlxwTJi+mqcwDU8ANs7Br+lPWE8s4crhDpy3zw6aZBiE
OL2hw1bJSBidt6JzoEDv0HuiDdNZvY9z9KRNtnayOxZaOvBwOPxdJdJJIxDQ5SsG
/GMYa5dZK2J0EY/r3L4S6fycJNmd678BAM+nKyYfUYPvu+mWeiMKwg5eMabKq59O
OKP/JTIFTajmGr5QlA5iNeJcKABxsB1nTP7D7x1kbTlQQsuGjHzv/HrTr25Mp9wE
btT1xk62yKGlatedVuZxAmWfjCf2xpKLk1PjxGQDlluF011CQuTtHFS2RpFP6Hze
q+QkbxROyAa1+3GNrgZ17fm2uNHAYi75UmEKyECYidpVAMMiNOxCQmG7BDxZgm9C
xzGj4f3H7GGng3dli1mKeAMwzVmeEOafk25+BebUzyyvrZ/fzmHu73miPV8nclYm
+xfnFGmN6jBlK/QQ64bDWrLgr0qCEOgC6rVA6+Ady68Avw8saAk7d1xU8eqybmAc
oe7c3eISMy7CZyWxmQQNKwFEPtjiKDpp+nzT6D+lyEVaBQFS797npKxv6D47HVBA
/zLWB2jiQYMuBAfCLQs+UfZoqov38wpKfZKrnAas9id+SBvDDX7gmgBzCBhtOxBE
R4ZUqjQP/QxaplKjL5UNngAaznVnrWY0VPIUC0y2/Tz1Jn5ivSO1mR5+PyMq+Ioo
dYbhdwn797vgsGH10Pk3AzY3ZWSPnqeZKBD4WAijPW5ea06EHewlUgitq1G4gMIj
sYhF3kbly+2IPZwJbuavd7IQf6AP+swJZdFJAEr0RnBkQp4xKeWJ21d1aLRlbeD9
g2Fa0x76U9AzIuWo0C3cEi7Fd2fq/pF6t5MN7Mlx1AgUpGe9TfxUltX1dQKR5eht
MfhQrKwu5UeZ/AQJm6VRyMYPjtJK+QorzHa0UiQDjB5tTwjjPAbm1RsY7rFxxpWt
7lsOQnFsEyw6C/F207zpnEKrDlWlHi7P4YBAKqC6r3yHHGP+Uq0LtJkpxGXM6BQE
MBiDNyjMu01vAy+xaHoLb61XTSQbIpn4wzyoJvfY1ZctbhQNGVJvtyzTlXgGvLTp
vLWwvyIUFwb4VdxKQsknsFwtqZKDeCbc0am5dyZBhnA5uHUq/3w0CX8VFDRF67PZ
/CXfNwuxe0ns22K9x+Q2cIOSiKCTqNIy5NJQiZ213tXgvdJ+fIREtTnXkgDL8eOQ
Iroig1d7pkmEXBnloplvFyjtxKM27FAxui2yvvkTfNq0XXzHWCNps5foN0HkNqiK
z10SN5CmKAfsjMOd+KV56JUO5cIujh0dGgRzhxppTt85/WNEcnDJuiIfdKmt3MUD
cIIpu5t63LtWFozIVuq5774XPP6LOwuPe19vjkheuxRtnV6iHXJgDzq1dxO7Mg7F
JGsNbEDwg8Csb0fhobSK9C+f+OeI69dHZp0uMNyMJ9dTWm71hrK0h23FaptSu7r3
v+WfmbBcm22CbSHDrCWPAsfD3Cs0cd0BQz49yraZ12XvGMom+529xqg0oYLpzfHy
bVm6K3sbe+qgQ50KdICLgc2Hq8fbfLr+qfGLrGVGnHd2r8vdEbBgj+SbXjqAdJUR
PfSuquwkza8GmAsSM+SxZ5V4wND454m/ZFFDpJOSYGXUkvFx+5y/4JaRJO9r5dLN
KuvPpuxVuT4yVK1yy+oUtRXfGEEQoFC64t4auM5pZ5il6wlyl0aBOHPWh45vVaDl
7inpNjIqY4TFEn9W5lRqefwhPcCkuJB8shSWKzFjsw6GknwxDx3hn3ENth5g/BQQ
X1UTVu/h4gvOwoWc75yeYl81U0JPklO7PmxBfLyU+8/LVyo+aArhdMhYxvTN2G7I
oWCBebn+rG0hYR9oXqDS02YngSXRNemV8oRB2219ShFxt8wlptgmk9KdwYfj/VAq
v/gQh4/1rxpfhFc5CTdxUDsEPSekVgUC4672tuXJzQ8TxpFoz7xDZAvwccKWlF9+
NLDI6Yc8c0HhTg123aSKt7IL6dh8whlyRxtskMSWOllw9jJzTX9jNZCkXl+ZyIHu
no7n63xC6xgiVNPDhUmX97ty9bqiQz4wXWxJRGcxVGgceZqtqs0DrJ5e3+BbTOF5
RONmo9/3d2qzj3t3Ls1cFa85M9vlUSJT6Te8lUPr2n3r02EVjceziePDAKRMcRUx
SaV+hxoakiPp9Z680rqm/2t++IYsMAiTSf7/ZTSDI4d98olBc6j7FxAM0qbHAjLO
1bC43fgkkry8aRjIrCfP2g8bm4gQoo6J7ONRGFO4+smlvWmUA6a7IqLdYkcre5ME
IDoyi27CRPaMnmuAP8JOk+T1rpQiQ0PCyGxxgwecAwDSVpo36o32dqG21JBY+yhm
jdaN/7V134/Tk6gdF5t0SWuGnOgi40HWnBkOjTQONdI7QnZZe19GeO5zij0lFJI0
VgmN/HKHMMjAjjy/Evn1EjEwxxDXieAQViD7BTpW+AVYBpKavi67WfCQbcBvn7bB
VHOfHLpJx/jgYevDb6y27EvOa14lKUEry+D4p9VIPp04nQdQZjhrkJ8eThclwQVm
BVkNFoxO/eh5SaaX/MeK7Kw0WpCe/GzoWEAK9X+oC+3H/o4rGmUYOU2GSXf6zPw8
Ayf5xv4bMT5eE8Hcr1xkAdM6kE7kqWa/yGapX5CkWHygEywcSWz471XNMDUkf7WT
Bw3pd0SqtymxJDR3zPusZ7Y0FuulQQWbI0oUDaAzHyvu3N32SbzqiKNWwXhZXWtp
y1dYR0MbpsVik4h08IwzyATUQWWimKiKaHA7TWU43iSshHmL+JoXLPOKsOx3BCnu
7ZdQeIgZ3Mx8+orf4NT2Qz6UWIoK90O/6Jz757QKaJRXCTzOIZuGlA321fHpyz0H
S3fSrDJw06lUBgCRYiJ/e9lE/4qhurhaYULdJ6k3+QFNcPIT1w9qCe5bHF7u5/16
81fIxGG4YJV6rB6EVT+clqQy28aFxtIYaIWTFihCbr/R0RrcJ4F7nDdQlGxD59YH
m5nWLNlJ65PSpA9TQ1dTfG7Os7EJ3OPCcNPvyyM9Al5qBd/D1R46Vhtzt4cCdkK8
1sbtl9Q1e7GXCqM2lhVoTFAYc6sRhE4Yf9B+SGhPe7Oj6dyfea2REuaCcwtMjM2w
s4oFWpM2gXD+nBm+eaR9RAzQS7OkoWhPkqT3+f5Fm0dBd87USFlQVTRIt7arO0ii
fZpjP9EB83dwrpsEp/umMD8pXKWno+tBs0HZP2YoFzlm6YiX5Pfx0OFefaflUyV3
RU/+WwsHsvN8CoTTEDfwa7w4/nQqm87E+GYt5WPVkBJxHyGddDISy0pbV0H+1BcJ
C7YlC8o1iyPgsv/XXlZS4QH+xMCMmczamMSZnGItuUT9903ktzCoSdBDN9TXS3Fa
KkuomnLiQeZf4MPpt8S4TJjorZBQpnjASU3PgV58mHqxgT7kTWJtbV6cC3au4nq+
hggGY8BVohCu6sXuAanvZkhgm6SRZHE1YMzoFVsGd3bOtTvFRRMJsP33jJN7Xmin
ZLVNlHFjPWmKWX5dx4ns+qiRItscdJYywv9Hr1/yVpMrdRDd8Nfcr8anxszwdOOm
PVs2s51rzuQFQW1623uYcekq+qb64M4CAFutBB4YRF06iZgCsBtlTwzIlptnQViY
0Lg+2YH+7mq0F/wW28X9HCSWg+BvktcbQK6fQpVuEfAzyCzCcgNtjOm/IdkHybwT
4X+THlClyGyaDNmFLbC7Yaaa/NNFo5wC+rsKY844trdmzI88oD3wvUdnMf5bZsRd
L9cdCfZ9Qw3Zal7QVPm6J0+V1sgmbUsW6MpdpOluaYYytN2fZJKAGXe5wBwWtZkk
DDBgEQYOx66JnkyTVtvLoUKpYY7wIHIVUF7oyxxwZ9vp3lXtC0ISxXbQXijXxFDG
kvuhl8Ua3ERLp3plBbxICKcvJrbP9DfzrOlCv4Ma7b15Qr2GWoPER8UmxJBBPyDa
g3SvxWfoN/rt9YwPGh69Nbgqsj3ziQE0Kx0WbVW9ao7Nk1He/rNRSw4kDFlR0sAh
6CwC4hyOYfSNmFwcU3KzASx379tt564IBbU5jNS0lE9bBx7N320x1AmSVvfj6CZq
Ox6xP0IAbnH8fXPJrj0GtxEOq3OGJ0Kn5AtvE9e9UjE7xEYPiCrJWQd10i+ZVCBY
Y8p35a1FpYAe3rp/3uXh/gEF8r44yWfIe5NskE+4OTokjWcVoTwo5K8rR+rux04k
cdolh0ZUqPPBTIHAiGvWgybUTYOQ4neE1dTXwt2/EYpxSXzL/MifIViayn/FwiNY
KPiGcuJh0wnmFe1aEpkTO7x308FeDbQnFXCchezgoee8zMirOtAV4xDenZYZeM0V
fiJHAEyP4z7Yfc/MJ/xsw+r8gfjjlkDa1zdpkqnknGH7cuKvU7v/jFD0jGAP7Fgy
q2K8IHCGEQ/5+xykxS0NCb5H++2LQte6+OpCtngEyrQPb0iuppJ7LKvE1M607hvF
dlCatq3QfZB57+l6wjTgwWA7Ks3pkBDp5PkD2eLygSbjl7M8exsdJ+d7r/b7n4bl
SSv0aQGSO3+zKAsLqcuw3XQt8NzEaXEG2hX4SlA+rntJMAXiD22bG84qlTM6owU5
cqYy16BCh44nChxXpPIrlfXL5ZX+m8uT5BHjiQ/SbJ+jGGOP5TYz1tONnh2pwWsy
LPj/mznCT6uvanZ7e7SNALPOqrKPD+IhIHFaV3UiaYlRVb33KNY60SwShAvGTlHE
QjvHLW7Zy/zGNL5pLiYk6JG9KZSi32jRyCPskv050jmPHWjQ5Y0/CqbOWI3MrX1o
J/1bN3CdFgux30Vhh2I3Xk+FsRuNjtmKg4VCzNGYvnxP9fe0TSNi6ZtEHpiWGbDJ
6jpegO79IpPspQVripwlhnWQQE9gydZvNTg/QmheDEgCA07BSQTLBZPvIrN0zuwU
Pem1DQ6a4mmSdKsKmWX8SqOP7v9mJywwzcoxh9SMHdvTzcNA2SpFP6KnBQFT38G+
zbbp8+eWDLRBSCXu1J2/t0zKSCin8FaQr2iyvKmAPIXSnSWQuL5+EW69KUWZnuEh
Wuiyv4M342pccM5H/gxMkl7QkRnmeD9a09A3BCTZNdPH8CHpSofnlALebUllAyYW
DJTChLUzDQKPEtVff4qVau/4c5xEfDK5pfvCg5lu5q3s3+oxXVZ7ZZGynyNbjf8A
VzUuZG2rI0UErpDkUCfZjG/vh4wr/5zzLQ2WoBXN4vTzqnzWL3kdkT/8TdpdCDQO
LKjHyRFEz06ImMizkyPgHM1MUMyRPZycogj93Md1jnYNVBTVTAbk1tDITTdP+KtA
8jqKY3MMcMMpaqC0pqgsqblRYXjG8M8BaWFlhVg5PwaukboMxuTUv/E7upXDH4Ld
4D4iiaL9YeOIE8zoXnOpwbNqv/EZGcknjpX2pg2dYJvAI9sZpbB2MuUS+ElXwpm/
fOSUuowtD0Z+mPgJECrLFdMB9N4HFuHppktzBdaWvt2Q7OLKtA4HP3QjgzvGBU5+
I7dHuR9PJpn/4OsttLG6qip6p6080h/m7wul4gOihFN4olY5g3tTsgVd++tx+8a3
69+DWjkalGsA9WAGk8H24BoImdFf9xIda6E82STqTp72lYiPEoyjRmOdaNGkxPBX
TpY2EB8GHI2sC5WlKBgmHjOfPMnbtXqayFjAXyqylEHrAV7zshcVsK3gkmUBBnNz
E3xkcwZ9vJN/W+VH4wTqNWzBVcPp6ReWF3msCq4I9UpeWHOeRB8gK47Tj2p3s9Fm
FcB+R0y/fmgV3auddrQFoFpsMQ1s+MnW+Uz/qTodvTUAaV7hdyh9w0SdXSjI+M2U
g0INrxdCPUxeXOF0yPxoTHHN/vrnuHx2z5duU5YYyNJiTPD0WMrjMjFu9IDDPn1B
PhHIA23LUXEx+di7kKpp9+NZMJlJwvirKTDcscfR2JKQk7gRqQ9Gl/pRJaFAJBo9
6ZjRFenNg+zRjy3zVX21w0seFjiSzOy/DKWlZWC2d+u6/CB7cMjxhndGudfr84b8
fmLgf1938TeGzEF8L/2fTCtCq314uFIXPF30tPtwMSZLkdFpbqzT3uOA/n50x3qu
iXryLgi79n9iW5rcxTyWc3xn6M38Hw4tyw/fqRjbAbo3lZB8neHXTU5NxoNp/3CI
9XJqtlP9rVg/IFemc5elhnGpBXopaP9OThEFaf69iz+31UDpdItuqOwvvPjzbXNU
m41xUo3LUtDwydPqyf2rCSz7tGv9vpmYB+/TmXo6k3MxiaBEVb/wPicWkgCJ79iQ
SV/vdTNItMNT1una2vAEJWUEefH/aekbcit/hwLIdFo/1WsB0j+z0/GsyUAm5GSX
5C6Ojb4ABh3nY3C1rUlRDd8q2K7ILQW39BfZu63wqOw21sTobE9fOEsZ3VIOimEQ
rUWVUxDAlre2Kn6mw5LUSlCQ9EzHxMMATiM47ciP5O+NHoGq2f96RjAVqwLV7liz
Ibm3kLBE0l6jEVPCCy8WZPOHCZkncnKgmVUQkaeXEdtKb69bj7jiAawWrGmRpEj+
C7C+3+xFgUIQlkfLxIEQjdaTZziEdRYOIrygwpwQGWHfgyCH5Hz53QWqGx0wcnU2
aetaID3BRuAKNbRDJYqQoOZ7NsONxJpIdQAhvjeNj7ODOMT8DYVOMmom35KKyqsN
K5UMteCxPGdBobELgQlT1lpCbK1cEp1uvkRqD0+NaNAAX5cLeEEiZ1D+RbcLxIrN
wVs6MCtxSOjqttOlgH39+4nWnHn0DpEZWSksbaLCWbi6LyjxUdCRAM1Tu6IsIHZI
vCK2NaJzg76acf1T7sbhit7hxzPk/thfyQIZQMh6ajo5mLpN/ZPtXaQXCbN9Jx5v
xzLX1aPv/ietGls8bSHt333lpCCb/JKBX9xij/QIb0S5yPtg/nIcEBbfRtKvK7Mi
0IE4EDiGbU+AJp838UqO7/1xB1HacIFE7+mYYXxnX3qySRVme2cMV1M1zs1oBGPj
hH05qm4c8MEN9F6NAX9hqS9E1ikwTByyJU5NPLr6n9mssPuF0KRrTsRc/a2OsvFf
3txzRPu8enzL/6AC248e/0Kq28/6nyFxXUDTlLTF6yu31zDvXSqHAiDBNeeg6GcX
HhU6zioS8+KKrkH8EV/fiQcjslsfJvXg6qZ4tDQEfWE47JmZ7zFJvw4Vio3lDvof
cu+nbRFW3b0HmbFvZPCBaawgMKavssPzDXt2OG1f5aDziI0kFOH1rcwaFnzcX3ei
/YIYwbFf8sAlOR8QIYrJo4K3IPbVWfuk7JIieht+RxkCfaB2KVv7uirqbaoVkoTk
wV1gPVkHFQH2lJZjzjAHVqLBLVPKmQ+bY0zuqFzDGSXCqsq4ANWqgL1tHzARvzbU
Ufzpd1qZEPuT0cImU8SXc0PYPu1KPc6RoJZog5V7SF/nfofPfiXnyHf0dhbIKJMv
vJavYOoHD3AzwiCj5OH1p7GpMDMAKk6HlvcSDQ4KPKWzzAZXtM65JrkYbJk5/Fmw
iWAQMAbyG7YbPPMcsyJQ39AjTmP3PdH/uc4t9XA4no0+iVQx7HfcmoFxRBNtl7Ro
oImF6CVDn0Bz+f+doYXR+e+ePXK8fU1FO/OBjQRBWPve7ZbayecyMkp6cszey0s7
iFwDv/upd0gzy7KIfsMPfKWn10HETNblz8qTOECogt3Q8qR0RDR40C8YwaeNo/AP
L3FmWjF1KlCKA0TAX7MQ9dFO493BJsm6VD2sh6iW76/dLHpqv9APH+EDmQ24MgfB
/YYGRBLDy4CUIH96KDshGKoezoHDnISFtTxDz8cxDdPJn6wYhB6tiN+D21cbIbWX
rPoEq21HjK9t6GgsIqvCnKkkQYYXKoe66pqHgHWBCjjr3JRh4PCV3WEyXPcqHcHt
w2p5yfkoVb0WYa+quOqOAnb1+GhL39qws1J7YP2/cWQC30B9qxL6SL9SxG/hpBU6
T1BTrNwhgrO9DzFC3UMhSz7ODGQlCTeMNETorFIaKRO3EqtLYj/7cScf0x0BFIfF
XvxyysRg8GwLJZ2EG01uWJ9ap1GPvLqfwM8VfW7SfWmI9kLoxIiCxTpw9DUzUOnH
gSPoieuc9VdiYoneHGEU2DrYU+CjdvUTJ64rwJB/09FReIDbE+5I/pB8YZGkyQ8h
u37G7T+At06NpBIi134Fg0XjYPrsp4nPm242yiHDi4lUjYustdrr8Jb6Iko0P4R7
7faa3sb05myMFjWk3k1Y0zYFGlLloQc6oKbJYcOFWB9VH0bn7t9r3oxjmUxjQYXM
zgPhuB8Jj+Pps9yiatB5Bbal/4QLBH35gs62Nhk8E4WvetgSKOUb+OmIlZMIFzs1
39Sgg5OcrnujfdnqTSTZSFYR477ux6nVNalbvMUEITk6Rk38WgB+QVtbqkD2l2Ol
aQyx/KD+1cqEnuqJapbuxhItOoM2lyeqiVLCanBfwYwcGzoLj/0+nAtWdhrtk1cw
iNw7HAz7vYewSu5Cp2aO0Pj8ccYW3GGjXVN5Phh0InilqkWhuNgPMMxAtjFTRyAr
JH0bQhNQ2NnrHDDEp4PHXzWwof4DKld/+SXBPvHgeaupDHoZYkPP3uwoyLAh7XfV
JrzKJ9hqGBmRGgLiQtr4yX51iFX+P3hzvXFpRgrfccpuGgkDDM2I1PtmJjhu/KVA
nuiwULwXYom9G6zWXNiFzWwhZW5wTPSOpqNfgpxoPD7vL+bwHceE7tvDzNh43lxx
w9D/osR70h6vMTd6KlQQi0WxNqlhDalM3opjPLVPsdO6ymY3FLIvPmx0nXrymUuX
qW/geE3KMmoLzrBcTp/f/Eco/adEJgl/8izHhWdLXfHONMuKlzttwyrLOHDkX6Jf
P/HR0CJEAHX6zzYoiX1rVs1PiMYplckMIrQfYUXwn7SNnlihHDtT+vqdr0ttgx5o
r1uuReGyEC78u9ILsbzOkqTnKonWu+Gpo87p0G0O4VIWXFObeeKxd7AyyZognnQP
tf28US1gUX+YxyyykVvY439N9Hx46xN8OSQC3X849KH2oajQMsjEzEOPxTl57mND
IY30ghYirhW3Rl0G41yyxI4HtA9G5o5HCAt1hgYH9GvjttgqCSbBYhmGSVELPWYG
VdlbmzF+gDuIe7Ute48Xa0xnIINUxhqJnO7QRc15b4qoA4iVgPvorfxX9/Ymah1C
+oydaQZdP/LWomKtAixRYhmhQqVMDOzSRbqCds86Jsb1vWzQ5tBDRSpoANc0wCOl
AnGxkLCWODv1iNrVvf9wVR4T0GG6YNbNsij4FzHtcUI+7U1sbz4B4h8itLCZ7MDw
HtGkD6O539YVZ3trEkB/M0uMoFH+0zhW5ptxhOzm03hyMQ7P4bg0aQp/2LmcK8wU
L9qpszRzDRh1iWUCmA1f4gRXq3cvzhGXaJv9eAPQEOb1JrHOH4YIKfV4QH7KmFHG
a9QpdPruS0yhJ5qWYrTGRiO6zzEa0Zk3gywWGdhZhStb936KDTTBsPMpnGLDKjgo
jj6psofHdKbZ21Cl6mXwX3VhePvmLl3KL93f2mlpz/KHJrKTSRmfL2ilK0ryhSm3
6/JdpES9Jt4hMkzkAfA08O2CjCYVNVBuUy+HKD+tm7kaZ3q2KlXWP03+2NkCzq4N
QoQwoXwE1GhY8c7+JBBFJsfeQJDU6fLVpGxP0qsflid3OwEqGMY6JpzHjtvTs/NO
CKqupa9Lux4HeKz4Od0FUPgEq8L89ZL62IUYURXXaLoxKAV+Vf+PUjQ+SHPtoBye
aifDS+9z2u6JtloSJTqmTSJVLThP42hMPbzqqhgDXw/1f4vRynxQrgiapdNMjEjw
9qKFQXctSTpdQxAZjWM9iS0E2Fx2HajLnvE6mV5Drtdb6MGdXOIdHYvQQw4oNkKf
afzgqWoLtCRLSJeHdJdg1JTA2KadnzL7KXItDPCBD6uakBj/daSQrGtS3V105Twe
G0O0lVmXklYCewBEaWTNIY61Z1wum8r1sja0ujpJEHBt3BwscWZJOWV8xehhoJ8h
ANJDamgPtFbGyKeotjk0qP7xyO2tDV8o0Yv+4zbSStJ+tBWHvtisczOoqY84+Mdi
Toqc5/1wl2Eg7CKsE25QW1LCN6vCqN2z2+8yLyhIkTVsNGUZBeYNU1KC3/0Fvnez
ELz/ky8dmfRJmwnd0p8JpHBroARNItMHUn1NSstHKoVQPelirC8bS4Whdno2HMEI
XYuWbreiNC1FPQK//HnQ2n0nU0WkDFtM85CR/xdAPRJg7/B7dQp8tJhi1Kvuil0l
iBsbn4u+mjmtjlpG+J+69TNMdCJ6F5Gk4lTbvQ5rfizPTM+6xlKXOszjNdeudA4H
EOvFhyhX7dZsr+cvt2l6OjdROwCPBbCdqf+MfZPUSF9PXh05hztPh09D/oRyNXCV
Y3oI8Sq9Tdy70+t6KCKIAZVALRFpqCEXgvhgCaZ2JZgJMN6E/9vm4WIEVWNg7x3Z
OpmUurlUgxJU4meN7yp3A5EVxmMFAXMT/G0SDTuZgD9n6xaqUd/cm2g/Cdl/s2Fz
IZLy0G9+Gv3MzfJ1hT8yBgNyeBitbN7vP0qGX+cRe46kdMW+15O3mDuCiSBTrGUe
1IE3Y3+nNwBCZCVt335dUO3v/rD08+IwTszDbT5TXKv80FC5ojxPHP+u3zegfvc2
mtEz5qNss8ySHJAgGLmexS80A8IfmMEIl3b6dMOoP2JBAvfmtlugrykq1YL+hvtv
2nEy1Svpl9rzLQIU+ilTv99FrT63ajV5u6cniS0iIJElPBYe8B5GiW+1AofRIaOC
JJr3eE3kLdTyOv8VJo2nvxppqZGvbhCB/gzkFp281BBzk31qJM0E9xEWxr/e9Wxp
RxN/O45xGC1JTDPdnwk3b+NmhKpiAOaIeIK/08KNyd9p1QHxnJeqovu3BRA4ZrLS
0DW0KB5Ba5tYIEfbM1oMhoiEnTSQSo8IPhArBHOhWaSq+yNkCsXIDa1XWsxPG2Jm
l+sUJbYmKxXuetWHABOprOP06riLq2aW+zsmBXXI8TQbEZr6ETTOZDTrYSRjRili
dvRjgivU9dCWhV/pawg+lImRm9o33gXvjfo/+Ai/lzEYjpU8yNJk5lBqptNwgXMM
nye1TiI7S0FYrnuNLvv89Cbkam9T8ZimtPd2EyS8seeBXfAwNbKgglTquTcVShZ1
yC8ay0HC+SIuPbJkLaaiEqpzhFsIQYBAKJkZR96COBdqJon5L1i/fL+qsYBsB+3i
Lc/1VdjxtE6D9RE9zgSVMg7IeCmtt6m/LRHCzTak10RabWlsethPSCZ2dUzpecUl
ZxxLRvn7WyKGi2tUSFPdOpJFtKROvFIcttLcamfSuD8guKIXdKRjHP2LAKMHH2A2
GGrI8xI+iH5y3XiovpDxzsSD6U/S5Rbg7lRRaUOq6LnHQ3l6L3biJ7hqV8NHDY6S
eqMrSRaN7lqXTVNbOIcCQ4MSlnkfNfd6QfJtZI0fw364qzF7cS0Dm1c5mI+FhbHM
vxlc1qG7TlEJZ7czM2SdKd0urCoTyGy+WSQ1YHOeYMoAHrJmmZrsl2AWtfNrJ8La
vhur9t0Xrh/iJuSwkedhkYBPShNReEhcGzHL394zUcuep4l9cGurgL2twjctUtJP
w78vJl3XB7j9lnfsLvAsZlc+KP7hIpKkK5DrZ9+ooUjTLsOXwK9U2U147NqRIIQt
zNa5NpB/4rXdyW+ELSu2MiZknlV/ZBpttbHmbpa8oz8FLiZwruo3J3QfI2GfZU4Z
8XwJYMa5NkLgyf7vvbvxxEDdQZg2UED8Bo8DKATBrv2OKpdvJDnW/w4ifi+lQfUg
0lAAlK7x1yIyAU8TSpK2IkJhsn8J4tfLYLJp7BarfJrqr3nxBlzKJoWgVb3cRNr0
E17uo1MxUi+9KIn+59rzupLer21Vc+6LjRdLFZ4OSTwGc2BprtJmhuXNeb7FQbBq
BDEW4YF2cepHdysAJY8P+51tSJkzd3tnZWZeGo83mq6nuaBpLHl0jlJ9jyp5MZlA
hkivBUPcnfSGkD7vjpWI2WCMyi9rpwwfiqp7PuQM2QmB6xrYaGLBJe4ImMv8iMEb
vtz+AevckhOej2ZAHX+OjN5EaVkrfc/MdfuHldH9I31enHDZL645zU5+lhk5x6iJ
iKb8/otD+yH/a/6YAPsvGTYEDwD1y+w+TGFoQl+S8BawKn4e4K4KR0lw0WXrYlb7
tWUAKMX8ncK4WtsJcKzgZAzkEM+7u1ideHKob0d+H3pdKM56NN8daB2IlU2lSySl
1uyyvwPJtkpsxqx1+22mV2PQqNLCcipe2Gv/NjNJ1hBfCF0J7ww4cN2oaIvcqZjV
csigx6IYEek/Xo1SIiEccX3JZowdhA93GTnmTaNUK21B5W02xDUcD+KJDUM3yM0j
/9s+Lw+Se1ddl8A3u76GTCdGtmmTMEu40vZzsEegLRKzJIkcCgfjpk2O7P1KteQD
9Sw7ov03/feTgdqZwkW0nCG66rLmtDjwpqXyGKPncYL9ObkfQybiHaKJPzL/Mxrv
FvbjfiyBFe+/QvQvy5uhgT03g+I/esDddj9SwkwFmGaLuaXBMmiusuuiL74W9wdV
3bCdH+cri0P8nU0UNPpWRrhE56YucVDAQGCRTgtM9tbA4vio3xs++h2ra7g7Oba8
jyYTxTCiu22ZVgWGNd3ht4AU9Me64AiyeYVxJ9E8WUH3X1VgvEItYdNZ2pvMtG3g
43+SAymCmP8uhXXH+8cfhWDLOKL/QTT49Tvdebm1Z+Niv40m+5uf6E16elWGS6so
y9yjTXk9cBkUxYc2q5vl9UoWvnsWdWDf4z6ryyRhx6GoS7MW69k9f8ScY6YE/ij8
P6rthColyX6aG+TkdlpFhvncQ6nee/JlAUQNrE21Bw0FSzr+jw1HwarUMOj7Ra6E
iURKZCnr8Uswz/34uAAMRTK6axm5cSezAh0kz0kWvx/qgVt5H7TfJS5hch7tfROZ
7nrN+JsH9FgJcbvxM1SGVYAaQYcI9ARM+/YjSRckvZDTqzZiyx+XEO71UnQ6zy+i
ws0TdDq3N+utvoOSFUtV/tCkYKw+kcx6y0sNAQqnX8neIIOhqySBr9wNj/U2R5vp
HbWV4Y9FBtcduIP9z0X89Ey6vJ9nuAqCBhCmk2WSxR63xhd3zykd6PAWuXz8Ytqc
2IK10vkLvGP0yW/RAxTxEsDTY0oFaO4jWcsoW+7XxmzqjP1ah3PFwc7/UVUk6ouq
evvh6FwoewNASuVhzWSMnKMh4PA+ZSSLMISfZPxtgfwc4bQXR9Idu/mWALQblTUY
oPO6Jo1Wrqm984Ca2U3g8E0mqoM3ORui5DFJh/EKs2hYRbDOGmZf03Z1RIKcYaNF
wmK+FZn8+yznUGF5vCsQCaG3pOiOAVHemQQZ7pFja95WD3El0dAjQvMBSRSYt+Ci
EY8JJZiJvcnOwMFmb9mYszpCnEQEJeuESNZOZ5p4ydQQIjMDjdux+6KiSwDsGcVR
ttmYwaAm4rjes1i3emS50lgUaQ2VDvhxHNrVtp6LazlDX62Bcgli9KlMz7Z09B7y
peWssC66lFQSNHVm8LXE+kvbHtWVIb6ZGujW5UEqaj53X/AvQe4Vfx3oV+Mn+HM6
GMnLNmAQhXDGgm/VMRCoHMDfOelTEkkr/Cvn4geZO4vpKdDBnDXIQQZhkOtMak9s
8gi950xxuHbFAklf2kyQOaxeZVO/77BKEF+RP+jJLtva2CV24d2abTVAiSurNwt2
sCU5ZF5tLRP34SNChR8kvZeSE2tAFC40w49nV2NVWrzBaAKmmFc4qCLHff2Y55eG
oA8DI4J7gGuMDkX+UMUgZD5Ye4fw3ak9T2qxifmbMqvK6T6YdFieuXSDelVfAJ4+
LZffsplMEZL/6jOeC1YGu2+a80qgwIwt204H14itw46jdSio4LGqnRO6PXmB0DY/
vMghuCjR5BqXmdt3OkGhwa6+CZUo/+/75sV2mFd9pkVg7qUbBKP3pRQtFajxRkuv
NKiahc1ax4VdsEIgq8FTb7llMY5uKHXE7+hpQOL7Xg27RDxZ215OFUZRLVo9nIGj
psR3Z/V+DFgEtmHXU/US8MSiJjgkne49g5m1ToV9Jrh6zloi5vXB0/iU2s+X63Uc
e7CWeNN+d0knIQksGaByT5E58312LfWHX4+lkxURXs7v7oH0CfUc0S8cTb4wBxon
PA1LRCHS762NErUwV4525XJ2pgGgastTxqz6rWXeB+j2niucvrRRdDOONI18k2sV
GznWQxy9dYXOhS/qeXRLVVhKItyzQthd/GEYMqpWAj93r3ZpzTGWuRDAT0OasE6n
Z+CQmm43lyHoPzWLqzypJKNg4KRunHZZiIKViumKAnaVzhwWfAX7rtVVI7xV/QSq
vNOrSvdczag+uwAYCXaiv280jzwWQ6PWsXHanSqubhkuEQYCgX2R2d/vHL9uX2W7
1N2dRwLa7058f7YOkce4iduyp/VXPHkNm5zWRoeEPcm5zTgb0/Ip7TvhD3OzNWjm
gbRCyad0gxmAelP66QgMW2LKbVRaZEvvZggBwH09HYYgk97UpiYy1MerB/eLCOhs
IlqtgbE2UQxgoifS2JmnJrGyaH6PzJKoeXp5VTssetAwkK5+7Z21O6B++tva9B0P
IdIH8Ie5B8dHt3J81D3MpYqCMCW5iTcLVSyTqS2eyuLk6NnTu6SbkZnHVlu5NcpV
EOv+e6UjVgAtgRqvvbT46bEYwTS9B/2iIs5SNve12Qku/CmuBiMFJhYqIG6+diQ4
LXxhgOFYso0oy6MKEvxHGY5HhIBWpV/xTtnCcbJbL3oqoviNg5YegcKjpMqVbAEA
MoqLfQw8uys1gbVXd4dcaGMX0OBbvK8v86pIlmcC4X5oR5ZYP5DNaH0y8SyI4VFA
clhdtzRLLtqRg7Wuj4pyjWO0hrbZMHifKGvYd8yZSz4fLXsZSLCORGFUHZPvmOEG
b1E3I3b+Dt6jwdUjXKsA7UJpH9sNIdod8znyd6RS2FmFyueHnrKOqnp8l9qFhpYX
40Oo2NwKEm8PBBZh8a/wV4emNdRCzned+6GJ9Uo88t0v5UcxI8mbLm7oXzk3JaOt
D2GG5ivl0CJBU3ey7VJ0gyzEh5HSjUtDOShGL7dNJDjF3nEQlIhEiw2vd+RfWeRR
L3fxxFrowrH4uPGCZKKpToJX1FqAB2dEl6ni9aEc8OwT4949r70/sk3UISAdpOTm
LEsRQTFp5tgkDKZ3XQSGTswOTjXnEwoSd8im37deUqm/D4BBlaM1tWZP0KTLHQ+L
VcYJ6nOK5rzYpBRLN8aKJHIKPZpq6hp1Vi8MR1LrxixJbW8pkLOgZQbZn7y9wml3
L+0eEdrFlfSTLbLQ7v9ma+hbDGuUKjs/evnp/w3TpEseUXmtTTHvRfI7OBTbowP6
bXz7bYp5x/4Dce89jaKH2wEeiPFcPnrQI1nHCl3gV8SQ2SCF9X0PO8pvRSLENlvP
mdms0kPoUo8I+B8ZMcGvbuuwUozc7K9OnoGt+dNCuuBCQBxGycyt0RZYCSA3yIvK
+FIZ7C3IA71eJ8PJdBlxvoSL+eCt8kHheBGr5/L6uFS408IkLMFTOOC8q56TRIZZ
CcQnKFnRfyF6NLZmxeOuUNBmt2QlYBtYLBmPYUeDqTy6LnTAVOU3paDS0pKaqquw
JrxQz8c5Hx0JpBd+AYzAv5SjFN0m7Lyhs6+jEzoBs6Utj71+ELBcIvw9woZr/mXp
Ly5oIo9A7v8iTZkea5KXMxMiPPzfMiu6ZajlweuZBNAqOBTOqIx9h3tgEz8n9W2h
sDaRUNUwuO/VUFuf6ezE5Dmcx+aOeHw3HbTXC/dt81oiik4Z1D/yXzoRhTnycNNh
22iLbiBv0Jzm6JKrqEYgxUSs6xY0vXfaw4Q8Yk3oBGi+oZdPY1MnrJbcciKSLnKH
6421IxUbiT8snpSxQX8UDXZNJY/Ju3911f1ywyxA6y3WNroArVCMFfR6sOJPXtFL
xw1f2XKPCzhtqdc5k1ojeVaPcs44uLjl1kUSZuBqtxeiBnRQlFxRBo/PUO7wKTzt
onaGkfBZKk1w6QHYExH7MCjQE123mp4QFuWjqrDsFxb8qlNk/ZDr+ww16+/3RrC0
oBq38ZogJj6GP0m8PLFOG7MS6h1CxDKrnodILBk79aQE00151DzTaeXiBwc84a/G
kq2ThZJUYICG+XzqaatWelbJfoySGhsCCPG5bgPHM/QPwTSPnNuA8ItuwZBk16Vh
GT7XXHTc37ncEw/hta6ts9oSXWwjc9whFWBouEblQrGAI1A01QLTabfIVQqVTEj5
ftKK4XeWg4rzssmpWUXiuItKIgyiha/CVUVOmzw1i3TPxrmUJh4A6I27DxEyPYLd
k/NVD9ZkGaTLJz9FhweJXOd1yiKy3O+vjIZ3Tyzic+v1yFxFWpyLhjSKHBR2i/0g
6kye73wjVgW1rHXVbjRa/LRzVe8OhHvXOe4/rUvVxCuy4VBJ1GEz59N53SKAY4bK
wETAvxwfVi2p4MdILYmSspxKFG27GMUQaFxp4a0vbgpi2xhEjakBXcHr+lp6xysf
Xv4EfQoGOTFCYZmhQawvI38z9guFJAIJX7uEdpUpKJFIAD7wBSh6uHYPSRmJ5gOE
C/45lKNCXTgMufY/GuUM3cuRkySlm23gKffWaOpavEMhmU2kE6BbitGscr3doohX
WNrd3HlzCyymkBges+1KUj3/Zvl0G0GR3SjWN2lbm+k5a09LweW/M/ExFuTUYIo1
wQv/IEvVpfrZ+TPm8UD/Eyr2LmP63h8U9cj0UtD+R0c6fNcepSaPtvfxU8hriZVN
rWOAIOzSBqVew0+hKk3a8yNVl5EHPDk0+QAHJsiQeFWjfVsPGzx70Qb3PI9bTgb3
S/cm/+hOcVtF+3oGKdLePA6QePiP0X/x+Cr8mP89o+7MXZ7f9KVYa3TxEOXRtMI8
FODzyBEX3M5KE0VLmy6+ng2ZeXkd2ZEjO06ObP72yJdBba0rKOdcnNO2Y69diTEx
JqcQgVjblA8QI5kKhuywxPXb5PT5znGw70G9lvNyKI1C1v2NIz1fTxgESP5QpPgH
7TawLiuORKDMlNwqIKD3p8OQ0/Hrz5h3xj7KLSb1PtTw9A736T4nvQv/d5QPIM5g
jQBJwpNQ/jVzHw3Yia6YrifDlF9mCxnJxUzFYdJbTHccVMb4Yg4KnQojZFzeXfBk
eJdJG1TIoha9dELOQCbIfdmSOtieUeosL9VukyLXKtdErY7YpuT0uQ6O5ZU6Z1/Y
71wqna1RcELCxM5N6njrvYqE8XJCQl1XNsEpK5bYICOhRtQEeQqXT26lpI0Uwg4o
0lXR1SsyBnaTPHCRadlTLbxHZESzssUMfb4FUvllg5MfAOBZAn1aB1GnlFWFJc3i
Q/xNN2lp+3/PLLiUjVkkZ1SmhWeVdfJa5X7JNSiBpeyZni56PUDHSAT5YuYyHB2a
9jcq+rv+X+2UFGEutXGWOxXtOmoQlEz3H1R+eFaRCOCTr1YzrSdvdVPQMnupn9Rk
F/ivwnNxPXtCgzd5yjW2VDqND6pE0m5UMY+rpEvIyVtpcmwBseC0hkcQRq6CU/C5
8CUCucM8L//e7pn7MRb/bxxRNftI3VqktNOO/D8OeMJiiKrd1naG4XGo40Vb6UIV
h6VuLFVgQvtKXV4PNf3xLJVNfB94zCptA8iiqMVs03shTecL9ycfjMAGrpihGAVf
3cesvFYbSy6A/Eqr1VdTnjs7NASTkM7a2dLJeqXpVUH5g2NjE6reogOo3D9c6MHJ
Xq3NsMs3jDMgLlzrUm7SEs0Ethv6ushcTKvqU1AgQ+BYml8XmTLBTWuh+vO6JmW/
VpD53vtQCyMcVWtFwcxV0OM/fvEN2Vm5fllIOOMgfp7v8YdeN820XozNkaD4fWeu
yilasjaYCGqfyZUIcBYAh7lm/LN0rRfapU981AEA1nva1PT9M3r4HOS1Jbnn+W9C
eiQpnxJEST0VmZReR3/Qg410jxEPr9HYpGzuMnsGrDhH22UEABZOuMBztXznm+f9
4gPhyQ6HM0p5c0lFgUocN3msvKT6bxbsG9JZ/78BqmEbAKVkowOeGHH10PxhT2x2
5Dm0cN/b+XUhxkcN9KnQarAiTplvus7oJM//wPgXdpqOgQjVvEya3/uhxg7KOAQo
P0rHe9QsWMY6wD7cp3rVF/k28VyWUQEHVlcJRmFDRLxNLq781/hag9H/fBBNsO7M
bKJh3VF9dwth+cZHgBZ4PpONTCRO0fZ8aENZJDDWHUJ1+RUlYA2Zy/GTZiawThOm
5Ev2xpLQHAqvfprw0Ss1sU5DUU2zlp2pk6qqPs9MiRxvZDfHIG4juqS6udxjBws6
paDEug55490lZ8+z7fTc0TiEvUWyYXovFtiBSwn9yePKkCUW3mmjVLs+tjTre8ST
s/gy3Zc5s/gQiB3FieLrcT089ps32kkTqHh61BNAbyO/nUNBfmfCdP7cIu+oFV1y
uW3FKsGz4rWyOdo2S60ShqpOAaqOMMgyNXchnaRxImoBJcaoS2xQ46DN+Si51X7/
oab5WanQ3FWUoEEoOctqgu4yx5NPJ1v1doX3sYIGB268UekmZr0/cLqlqnwY9ptG
ryPSnnf3csuQHgtQF3DU6364UWWG469S3jge0MD36gVga4kawk7kZcK5eeI6rbEj
+/Bc9Ar80W+PnwFCH6RKFXqd9Rn8sS9BY93w03PAwrXBemrr3pUeR+kzXaXck7Mn
9Ko/OPZAm9R0JbTVnQHG18U19o6Er6AGY6CMkaZWrzs9pQ+xmXGCIbG9RrbYPwRT
Ijqtw13y81maaIZu91FR4BjGgoNcD0r/m/s356zLGKbXD90TD/FFyFajDcybbHg6
0HpgRjhipjp3RFlD/uKdZ32yiiZmjqvOcSDMwA0AbsmuJR3C2HLLWQi/OZ/HgCTd
PbQmnFxlLGz8h7CtiHoCq00jkekYu9+dl3ZSgR12xBdgIY65oOP6/OWeUYul5qsK
fGZmmzrg2iFKWXrBNKyH7quBg3sUxITAUaKvsH/8p7NiVsKUFx5ZhK7HrolGGj7c
sOGMLKRBbC/8ZAfnnMfAPWGHwUKFU432HUnJUva4fXoR6RYGWaVPo7I0owQvn7pD
4IB0uaeBGEjmKVQqV/iypJ7UgwIFsecwLG3yhDaIme+4zLtIvr2VHyAE7Ed0OMpL
u0MYMUWi1+KPdUssxWjEpdhxC0inBG++trrwMkFCpwMUYQbAcJSm3ezRztipAduM
84cmhF9U/HVUqtk6d8n92DE+QTz+LfbsF4U+hR/IHkJOaKYyC27sbMoj4iykIing
4O+31PgE9jOs+PJ62C4C/WbO661PN4V+MYarvditoBO0TtTRVpruHSZT2i8GixJ3
79klsPNpvOSYXVOkP3gTkyRE15JnM+iDc2xs9f14IUtbAyIJQuFCPQrjOH8CBNAe
hwxT9JRWxTA2WNpdT5PikAemWfS3vySXuNU6IR9qma1t1V/ZR6K54WDTGcpY+tHd
4DN5vZP48f0fDwB3Rvz9dOAJoqARJVXqfZRKbdKoenWcMomb1lCTzWo1WfRg2gKs
D52FSsjexqY3S25WHI5Hep6lwmrEakAjmhQs0r4uLJ4GXS0YAz/YsxY4qJreFQZA
RmDfycEVsNFMkTd4yYhTonSbLLr2/nm8kVO4U3k89SZsBp+nvVwgqOX2PqdQCnrx
QwgsZ75eFVKZCmwDhgLlyVnnKX1T2Z7YcqsZAHxMerth9qoFONELBw0OFnwAa1G0
362O6h/c/PaiUxw0Ym31VNtbCXsK24A4eHwe91/ExEuSWJjKxhqwm5Hx36tj4jHr
wzhSlbsortM18wRvU0s1q9fXgvo+DuzcXM8iDtJkvcfy+MwCbOiGrAwVgmDMDCqY
yxJiiZ/Z/XCw77Tpxxp3soQMTU78PMtLAlulrPOEonbihclKKaYzbiaRzm3aG+LS
HwP5c+gyf9JDLWF2Rbn561m8maxTa6dtq+LulzgodxuexQVlHXuRZYQvVgzUygY/
GtvhOjSPap+ezSXo4/F57qW0pHPZM+pVqjikvk0YRnkDL5fw49rD88jFnDt3+q35
Bco0FrivZFIDiCgJjZFq4tVc+X7OGHPvDXoSEjjpsUGxMVuAjFMny4AYphYJ9M/e
MI2ygZqh7mErZ+ehwS1YnGp+owb10zg4Cn+JddL7vMFVqCP0rcZf4iqPvzQ9y/C0
cUq68R31CxLA8hZX7G+SMfpAk3kRMPUYlhwyODeVtq5kitu4OGf5+8GyZ5mURGtB
byUBxrUFv1fCPVsutyKOhImcla8/Xsb/N+QKaAOGRP7WrkRm+3PQPEyEXBMDkQ1L
aB2jgcH91dQPTT31lkGtAyNTYWITdME6u2Sh7h1kmN6vb8GL/7n33JP9EPCvtP43
SGsnGHVKlA5vbm1xcmm9q3pwAVubdnO9UuIxkgMJ7skCaZkA+jKbmh3mSutZ+nDg
S4mblOCIl2l7v1FWMXGSSemGCohRhGQfhVnVWNHK5jnSVuzMxo0jHgw/ekLwvddR
n67Yl+jnDJDrvyYUSU8TEpvzcUKmy7Bz2yhtoy9ahvVw1ETr5BXL144qMbAqHsGl
1mjXc3KsBNL+92AeGJ6NYeTSdzUNRWFsnDB8FFBBO/wg8Sa1oEXQRGXryR9iMaAg
+qnjcs1HG91OVb1VIQomonFZg849dKq73XsWIgU+G4nBB1BXCNby3noXTauS8blh
EWv3X+KRYwo4GEalR9GKAjG80cBuB6BITQb200brlHPfog8aR4Ok+7f6Ijz8Qt7L
IE1usbMRV0mSe3TMilTXyOrxyunmd7ZHsQ1xP01UrD5weGvz/c0y+5kf39KsCIqA
eT1UMnC4cRf7I0f+3Bsw0AJ05fIGphf/Vgkr8kW+bMk5vmGbhBOYayZg8l69Y9Q8
8VvYxuTGQUxrC3y+dUkNKmowR3khxFmFlyQ36uyPqp7UtPAqBztxFZUrV547reE3
av5OQzaasw8KZh1hvK0tSVst/khatj3+qy3FK4ffbN+MJHXg2zwBEjVmN9NBR+bN
ymE7An2eHYL9PKKcqK7tjRAxKEQuP4mjjyIfFb+JVSzcpcouLdbp/IQH0UZW7pfO
HHmrleLH4K46wPtc+vWZad66poP6HUWWkhKiU5hSBceRpPhYLZ9YEuM627R+wO9O
vivrTA+RvrsWxs3lsGfE5fV/2yrNx9mzrzlp7rUzQpkpJNI4QT7GcjS78xvbK0pB
tyZNHjmyQtnRdAOm0ba7CT26Ts15t19SvjkZnw14qE22jrKQRUYUZgYE15VchgC4
R4aXEIB55HkwTEEF/864c/CDjOEA5BEcPJ/0dhvCIQY8jYONVQkIEwyP5PD9Icuv
qLIAcnGOGzcvllsB+3+YHd/MEHEU5E10R/H2ed//vdJx82ZtmjksniC2oADYysMW
s0Jd0TtUPm2pMTl+DgWotxVowfHyqIy2Kd8IvnJI/SmDTUi8/Abt1pUURHfHF/Ar
iXoR5UOoDHhCrZfANXg/wDX7vWQ7pJUFlp0vHznC7RLctw0sP5Jv75u3e5VXu4Od
ToPiZjODGyhyS72U5KVEtwO49afC+sOmEbvQeRd6lgzvwWme7v5j3LES5zlruwNo
NsJmQA78aOFAl1Rx+1Q3mu0RxRkukTKkdgTBia9pmPtaumZKR8TAFxXTtHcedTaF
sX51DXDeJZ3VnMBXRjlyYRpEvmA+61F/zLMWcyzyYavzYSUATlgGUB9iwADGyh1C
Gx/bZtkdxl9JpmrJW0HX9ISZPb9e66nnZ3XYlm45xropuG8fxWXLXhFrG+ZU2RNq
BHXtJ1tlXmS65cfxV6IjxRmrvHH+bCxZXaT2/L2yAIcXKNZkRKzNxVKKob6WHBL3
WLq6qJZNslEm+GVzYKwZnWJFfcRKFNGuQSVZe4CH48/qI/4lMCioeyKKw0fzcl+h
pCZio62BmdAeLmoUR8L+J6lDYE2Jtk1c5WNp2q6HtNo5b3Xo4lioV1sf5eQOy7nf
Y5yK7xtHAyGuJ5uMqmE2KRMH1lJKZ1Q1ePrR/XQkG6e3/RT3+bONvSg7lzN+Eswu
l/Hz13q04RvQ6M8TIyouylseiWytov3zwc8ccTl9/iYvUnZ0QvQIByOz0rAM24J+
4ambVLjyfGRDJpC97FDaZhDNEoLd+p2ZOIrxsCU0xPPTdZ8/QRPh/iZpq4hd7DG1
PO72YtwBwxXXHoi1rVeOtgLfEnjk8yErTrEgXhLhMaI3mBrpEKRkx638Jgc1RkDk
P4kH5CFmVRNr+1mj8N4tNKFFHT4/M/T0WC9gJMwc1mZnydWZrsQ5t2r3u7BRmfx7
7WWGwEAScdTuXCiujjTfTLoMz1WIHMpFNGq9iOsZvitHmAB8k+RhggPqeTmzsnfd
3grvoKppWMqCtjNXuliiMoYfhEzremnRfc4DS+Y+i56BeBlSypNws797O3Cx/5en
08vgpVXLDfdrMNL24jsuib7P/ynQYUnCEaEi7S4Lcx2+GPe5RrZH6X7dj9Gf6Ddp
tmO1rV25kAyF3jHm+K4BxN+eDjQARTfCYgOpvkpfUJx7pspkIn1NmCMFZ/5c1dwb
vsJq07giziWDE4Q4FAKGrO0yZdkAaOrqLRHScqXunQod8hhr+8LTS3X4+uwqjerU
jGFyBFASb7gSyEhTY+gtUFNUBV3xw8PnPybs4iD6m7QW+SGBSxefZRfzfog4id4i
AZpvApa5Ojy0+0HrcDQtvgm4MJeSWzXfpBUlQ5pxPMUPOLr49H3hmUZjvI8NEqND
Y9q3WWABCfEulU2F97JPfItdPHARxysw8lNnF4W3H8Xb5YRd2ZfQ/0hB1wSByZVu
WQs8ZhIWZcJfrkZJWGGOZwnQ9TcndiybL9RDE9dq/iAZ2SxaeRCQPQtc1hyBfuvJ
9k6XjRoTcdkNypmvJd5KPNi/UsKGMHyWE4QXAGY9iatSGSvGYthkyS0JgxVjThXs
0C/JD5dF5JyAmQRQ1/cZgzlXZuP8fevH11E4gDAF+Q0JqY4bvzJHfvn9l2qMNnFc
ZvsquRGB3CPkW1Z1Ys566J6gIDJFAalwjz/rgfE6VBfmIe/YSllUcT8jmkK/cSfM
dzdiXLOAvePK8y/vsVILz17QC3tR/ky2omO8FFR8Givfyq6ZCap4qEqR8u2WSP3E
7w9858Xp/qQJF1pKGxF/PllJT61nTyezmImylC86mPN9DDr8MuLHr8HcqTqSQZoP
6w+VfFZcWVHCFgQJehYU8fXDGhcYhOaJinq1bsmBR/E6WU2xS+s0tOGvfq+wmGpA
o9df7F7UBLs0Ml7BJq1eEti6MRkx396YbV1WGwZFzhyebZ3nw0nQrpyj6NXT2Swb
rf+v4W5m2XO0sCuiX7ESJ7RytKjWWMUNct2i3BRGJqWHREEpFbTO0bzEiK+NDL0F
vtLc9OU21/zuO77JiYbudwDSSDpCGIs/KM98eIlNYMMciMxQHrfq1kQSGTyigze2
2wK7ucvVY3f5lu1ZTo/IBvgVdkOjG4h9piHy1O3M+7r6a/IYeqVFSPqyKxHdnkNJ
KnRM0Po8PgSajkKLuqxXpebusgkU4GpBB77bF+ihbFuap28spKr4ABWNJaFlzT0V
i4fkK+vA/WJ2uX62vAub4AR1h67G7cwopVd0S6H3459Bt8dGN8EXrz4vkj0wEgpE
Wpc3gY4w/1wLlbJ1Rb9Km7OlHXXzcegHkMlhivDgbVF5SDVnQ/EoJe5ewrbJ+aOJ
LL5OmrSAPOhdxtPfCMIf+y7fR8TGaso5XstmopiNcsQKTLsX7sH6EZsZAGmp4CBn
ua8+bxPzf/H+OChsv4gNgdno2dIgVPw6AC6lpwZAjUyHgnO8BUYZ2wjH3bmZzKtX
WNO4ueONkOMGFX+oRaWeGy3FlbYVwFRhToJgNPhATbrs/DEcLjjhQAShyikp6Oke
BepA6entrKZdeo++mFyq02IFmdr+dZd0gOWsSl9+1JYfc075HkC2RN/5wKCywwW1
amLlCfwufXSiKwy8Y+AzBPKe2odgo8V4sBsPFtq28EhLUbtjC/WK9PdsOd6nDtYO
doTFWxeSTMLmYnXwFhUdob+gMKw87ryGiiGGkcHTSaf3dviHxVeG0KD740RAgxQi
mHEOve99WCv2CFi5Qsa/M4ZEVxfs0g/PDQNGreI0CHQ3+DI/dGI9z8ywuRydxbH3
bB/fji7VRupevGICIZpw2Qx+JBhXuoLPFmFWxo26p1wn2Bje0+5FvfiFl26eeeFw
bQkU+bpKJBuTGRLmbLHocdmbTttHH/KiHlbkZSglvPRHMJsHaR/Vyp60CCQ/5NAo
ecnXeRRewbs9y6z59kSLPl6lde7CELOYBY26+v6bLAzqbkGVqXPaNSg0EULXpVgq
cNrYd2KMXxKjZM0fRLJZ/fqxlH+zBtkkWEGYZFpBvCR6J8fcNKA7jNJZVLcVWsr4
oLFsTxm/op7P26L7CyJNJ5ZwU4ZYWPFQ9BsnMCxEX3KS6FDQ4QxdZaYMAzMSK0Wn
BACouEojGeibpNaohJsrxwXsh1cOA4e7vMgh8oPoDZtAZ4ku5m0KvsfDs4g/6/rl
tYcN/hQaBhfsL499cOhZ6qwgEuNww7eU3sgSXGKPcF7E4LiEWmu72Qpgu9ST8IO/
ZN4IjEBvSGJv+MN3cT0XLMphEShdfB1hhiPVPOHn374wpIQOmXjtVWRv8p7NgMmS
mBUrUpzIF6oUe4JtXMzqkkRjBsgMIAxumvkLTGWjMZ7a+2GPWdwbUGxiPvmV6eRS
IP2fm31WyVMNwsdtPRZOJ+TqLHRvZrQP1+47xJIudb3EK8ZvdY/92LAsBYaagJP6
Ds/dNOq2qmlnCQBtMfmjMHdn3Ti3omufAgEsTMjyUeaBLQEMjutzL+aDErhJlemJ
Z+JKTS6xhZh+LX3eeyfanAmGRJUG7emkx3k5bk6x/FNeiLumJQJ06C+leppY2XWT
pfm9MexZh4Ad3WFc5n55Mqjah6ajck95WHmoHaPvWqV67YOq7pb41DwlZ8aIc0RL
sfiRtY9i3L8Xo6w96Y4ds0UrnBLNb6Kdesr9pbcJ9Y3shr6G1N/Ut661S6owDOxL
oBPXzhI5N01AqTymPaayNA8IFS+wX71spPehDVBj0nRgySDzhmJzogUqa4gq3akv
VaBhO0586OyusvJUCqqN+JEWmdAL8JV7h/Cav8dSVB1oShjj6qlrg97Rl8/o3hgB
fsHX3BiP/CWz576ptaJuRo1/XRCV50/L8IQPIJtyNaelm3oCxfRkKBr1N0LAswu/
j8zrTie+XktjCP3H7x7L9H3Ga35CFflQE5Y2ZYeMK7f7tvPycP3dTMwLbttIqK/C
8HdeNWr/tGoyoyK5iVOcQT11tEMjLx3ujMhlRRjOd5Foj+zp4WP+COhn7Exxh6x2
0YnJKhLabmNnqFdSQLUugD+m5EDZ8HxFD//pOAZkmxKy6oTB3zgtAdBdXbLXAr9J
nVYZ4uXlNtF23O/eVhW/D1rs2E8K7K/958CRAB8+OJxenOtZ+w9GOAuP9vBBlxQO
veoOO3pvD5Qr0pHC0/GoKp/GMfJ1muD5r/IrVnsWzJ4UEUmP1gcnLHwJcsgY9ZOc
kfuRa3gh5L83cIqqN3+QhbeRl/7BTYlzhfxRJBzjRLzHeytVSzZlQawy8VXLavGr
xCdYsrpr+BUilsnkj695c+x8JjUqqWN9cU488sbvy9yVryZqfrdEKh8pZj8Zkx8m
JdL4H56bX26AE/UwyC/e0/N4RzzSnyemzRZlGaWgiZDofx688oCDgzrdWkr5DwOg
3Rvp6mMbHOXlHHU1ZUcyurDh/WDTkL8hf2SzQgvjR75Piu7a01zPnCNN067YiwQ6
vuJWDplsV94vUmbgfNljStzEjAphElMqeDoAE/N/GpyAlrUMIIysV5zogvIqwtbm
QIzlQdn3hzWK9mQSj15vHUV+sMTnf68mWObNWTMIP2b25HdqRkOW8vlTVmVUjSWD
BtS1VdmHgJp4OKGYQ6dquannKCkUPzAVNLouR8aO3xhD4QGvcIq7WksnHdr6spXU
rgYi64pT36CVremzw2z+24NC1Mq9EL7AEWlf7R+/HpNUUi/TmsBwKNGJT7xco9bp
Vkia0lDyIeQfBq2W2BCHWGxYzsYNbjOmtI+QJ6ICprpxSkhVgN2pa++Njqzy5xRI
xTS1OewiPYcTrUTTZ+B64cE14IE0q3FbLlTSFBgTtfrssad4nvqFSHg+kkn+r3ch
xRUYzq8ERuwRRR17aTcyri5gTP+lyRfvVsRr8t8R/wEW519kSej4jLGmIHE3nglx
B63JTTasR6kQy/F7zNxXVIZIRDb9D6GAI5o7rU068qCMgglFquxMp9AQMhcg5DG3
571hdKUcq1EDfJ6gsOLYm+a+LC/MuL83zpLmaLawXwkdrmXLParLHGv2MS8XT6ng
pOcgbSyd38uAtgqi0xApdpwsykAL51gfxPMLWDSZCn0D2WvXbWy3YMQsk5zULKXX
kW0uudrKsVrPNrCbspgTBj3qc2GNRDEvFxie870W9pjWhrn+UcJo5ayMtFJe5sFR
pXWRcHfP1RTlpbe3O6tCfOx5lD4gE6vTkYgd2ZykjU3ui3GaZsOFt7BsRfXMp5ak
gax4+NdXP8+vw7FZ4Hc+UOpLshYLf2B+H+DODjb7kspx/1D5GX1KouIlFp0xFLCS
jT/BP9ZVMPmfvxTlqnyYWp6//e78SFFT915uwT1+21lwQUj9WaXVZsrKM31UTZx4
SAMV6w0NVmEyOp6lnBEQ6MNehuszvf4pKtKKhp1XkTKW9N99Va5DVzqKjXE9yIig
ehjuAtiWxM31Os1lIChrUn3YDfKA0k29YkY7k3y/PbWjEH2Xi7EVeArNPUVRPwVL
zBSYFoYQ9lr8veL4VLt1oGsawOdknXb7s5Fmfheiie2fLEDwV9EcV6/uwEALezVc
pFWsLS9bPTCrFuc64ifhSnxkaNwSB4L3s5Wzu/Ca+xfGoNQuL4Ely2beYpqHxw5M
mQyAXSMmakrWrzGymKLSk7VdESGp9yRnSY4XEjq/5lsHCArGxSNhfjKuuF03ksCs
zuXWKMMdwA5KKGw703uO7klJddaOlcYu+FcGtz5rIPc6PrMc7RXwapW6uFOJGIgB
OgHiYzhADFvEb45CqFFpvtN94NgqkWqhFUdpEgZz230NpcWjcXR5oRiSAPCJ5m1N
Td4Hir1v6nQs+uIg95lFDEW3R06xLS3QEb6JBbZDbNF4TvbVFTRmcJIGTVwtdkAk
IEwUIGsYtMWhk6EYjg6NO8fLk3Sg0/I5AfMnKNW1rgeTFg/Ca4mBDD1Y2b4o0BtN
Tpe91qHeq2yNoAwEY/k9zJWceJs8OQjtpHsJ7TJFbA1yRkOd9v2ApTdtnmBOu8CY
wwKaO/FZS6m2uQ5zWk9omJncNJyThfFNCiKJY0DsfQEFyCcbFwuVwEnvgQupQb7l
XnYkPNs+jSyQQgVPncymR/mW9wm2pTGwY6xqmZaVbs1okK/svkZnoAyd9yhae6V4
GBoCU8PKTgW5SClOkJjK48AUdi6oiC2qq9wOvQA3gkoe04nkkos7w6+mp+iC0cML
JZTfasAE1R+YJJ7r/Dvgs4bgyeXMsr5ZJKU/HSRxxhwMTyE7jpD4xE9R1NMZoiHZ
Kc2NHG8jONTjG8ePUeUH+JoDGQ4K9jIl9OehoLCmg70uZQLL/1eh5G+7cdroAYq5
JbkhtS8mktbd6sYVD0YBsv/Q9O9/3nrS/itKfZl/UQbBT70CRRsdg8Wdpm1vBoEi
syAMoshobre0Z1f7M6s65E0wCli+WxbrGv0kGZtE/6H/dF9Nh7qoyrV71ieX4u5/
YlmkG/GgIXEAawIJmUVoVZ1s9k+4USFsot25gwnHzyvrEuQzUxtyn5BMxqcIoPdY
CmUlzqXf1aW4AolEfHQIHt3q+Z+UMDqnj/bZ7nsgX2RF5qwjwfybQhEWGXKBwPWP
RoqSOmqeH5QeKdoX8bpTWs29p/Ipy5ynMwPBfrkCBRO3CY6eipal1W+aXrhyUXx2
86wu34wHkcegSpbDfwggUb5FmcHmLDw+AVekV9oWGqUEeUdIbqCLNEauAzUgS2zO
LohruCJ5OuNXnDWzxNuJxQJzgyxeFFOPBjEUnpgyVQH2Am8tEuhT2ziv6edrWd4I
xa+xoifUfzIDOAWviWc2tZt6AwaByqoRAq/zG+jeG6fb2WZONn+lLQsBNUpbpVif
tE+FN9iPRznoVapsdtSrX+byfenV2NwI6dPIHDt4qey3cW/eBpWnu/4IWwiLozi4
Glt85VANO5z+w1cmGHxEoF19ZdbrbgnsBz6+3PnN1lGPmY6NO8EzaKUWhLXpS5my
lEr5hjxuSGdY4+JI/kSsOFC885KF3RuEiO6Qq5YL/7Fp7hsWwMLjp7ZbKG8uClKe
jnAA2ZOJUiETeQ9xndMswkevjhCl3mZC7ShlsVK0B3sx3yQLRBULekvhH2AshdLL
f5tYoX+AlwA9gSmjs3c+5P5Rhrj7fyx9Tqey57ahFHlhu7FFOyW+wZTFZs7TarWi
tWGdG9cj+x0cke/7lYUIXrG8dAY3QgvLbbemU/a86MBXsWe7UcQ7rbJ53+5KIVi6
GfwBv7zgnn86StQ7zkteewRSBbw67i+Hmc9aldjxBGqGbaTLV5bS093DSf1UhEr0
ibfnF1sGgeBaVLHJ2Y4BYaFRQJy0r4b/4WVwPDjsRLqvRlmK+ui4o2jXREQQHtqF
Eyaxx1Jpp+mAksW6IydKvp33WXoLwTPrE5OD8X8P98cGSJtROErH8rjjtpYi9NHm
ZRsMGRnSCOYF0rTpiU1kgmYppLLViP/t31lJ/kfQbigE6iTGAfv6OstNIOe7jYTB
J58sydbnplBX9z6v+yTtHMzqB2JIBbdJcARQjC5limhSZWolnKvp8KrlEZAIVXUE
qWogPKd1DTU/hXAMDmyosIeZNScD9yBrlOiKEqoOanN+qrfr8phYJ+SyAJ20p5kk
n1vtF1XZDhDS/xB2QUVXq/gH8AnR4DVM90PdPPH2OteI+BPWh9CtaOVHUHTGMxf7
D1RKtXzhvBGJIjonj/4IbKfgdgB4Ke6vWpHnSRKVU2ZQvQ4j92GySNKH4A+Qh473
vQXmxJs/HLSUCg+S4jRpGfCKHefZAucc9ryC16VSHu8ZWqY11igYAtPahoJM4qOR
18/nYw++brtdHGyBqsNZYb5HWY3W0KVwZEB4QF1Gr05TyQMrY5mSKsJ+h7aFuvsF
ke7pDyxMitY4fVJcvjftUEZAf7GaAs7OmjGYREmTscCrN0iRCygJoUeaAlfU/ln4
Febr0B7biWPQWklMRh1aqtgq2Kw+i8Rom6CYfDYeEr+EsYXJxWKhuUxTuGcRRhrx
+Bm4+zMTlHYl7jEaKD1WxcWggn6VGxkacl90zzdzP4WTY8b/+6YwyduZF6b2D4ao
+qN97IvZ90khTAyawj9bWzf70/ZUEvnWngNpiJ5FdCyWuUY5TgBN05LJfY2lmTRS
JBgM8Lky29aRrfDElmhRgJ4+QIsyh/ibOu6N2rvqzfw5Kn3y3UQWacO9OrIeMLgr
inSqn/hYNyQCczAQeRgTTczh8iZfw+2VUIJAxy9z1+oylL0PAlspB+kjtOrxQ3S0
+z5P8EY3hMeA9MW+TfLXpjsSDsAIGbQblIEcM2hlQ2S4FnRejOPz+aVG7ZCzwJDO
BgJ01c4cmSGyW4jVLscSvcIvtdhwBHFy0qYSC2EnHNaXjCir0mxFzhUbXGcp5Wnu
lbWRl5iWftnaglrj/UxD/htL/gbAtVSPRjvFGmxRhWC8zZuWxoCxXm5AWv+vy3k1
1lq9WWRTyfqmTr4QG7yn/tpImhwRj+Lt11d0Gfne8sHip24beRIOs3gjc68BAftT
XFIpAWLknyba9JqaV9GXfy58BiO96dQWfsqhB9Tka/6ayG2W8UPFhzUNk6limknP
7ejVjitXhO/SvtJCoE2HHeJK1eFo4RnkAwXlaplvl1TOX7UMB6Cc7NOxtYn5ZZ5i
VK5bI/2a0IBBm5e90W4JBy7v5Q3LPATwOc8lFf1HE0HFaEKcZkCqnRMFhqChxt9Z
xnqM1C4PBwfcNCs8jbcFJ/cHuGCnbv76Zxk+ftPqTe3pjyXoB6x+yrS+x1GixOlM
tudMPAXyiPF1uT9/XrTzPCecBDasjKPqCTwI1y9WrUpg0N7+O1BP3CcPvn247Tn4
8YBnU7Gne5bB2Dyc4UC74xsYoZ0JFTx7fUerq99Mg8dwH0oS+dIwmDNn317WTKVI
vY/lpuvcSdJIi19DlAz8Y90PZQiOSH88kAAL8Y9Z10RVZ0Gv1Ovky74FqbiJF8ta
hv5lUUrVvyEgkAH3jgkB2Aa1XYY/Exn0CV8wW7YLZQ7kb0l8Qe2CFl5hHCAVcrWg
TBQvXZAzeXK8ZgeJU6WLmMArScr7bPyuuNc1/rfYQLTUy/x6HwR9dPt3/NBmpukZ
q9gW4FydY/HLtY0xpGRWhC71I4dn4e9amHXs5rLWn36Zs0AVJQ0QB9jlrnBq6ntw
9isXduLYRbUaQ79lyy33QaNAwbx/goRhSmsJxXi+xoErxH2eXfGAGfbfymQ/sgLe
eXXukZmX8nSsSmW1fXc/BGB/D3F07AH5Crx8+cfJAzAntGiwGFsLrRC8M/0DBwk6
eR26nRoCQzLB6Ha9cletTIpAZ+cpcfWAfv3aNSpb7JnGtHtOUBsyan8LkLXDRQW3
vnJOJD8+9tW+7jdugaxGSVofsfeRMcdfGvoLlTUgAXuSiUbum9TIDTvfhaziGxt4
Al4JEN1L0wOchs1dJyFWMuKfkrHRSJQggpHcvXE4dcDLf3w4JEKbJl/nJXgRsV4U
ezfmLadYhP14RNP2ki7pSC7/B93vzGg2g5V+4qRAVjg8dSPngxbAH3EH2bo2WeyK
5sFaiIQhLqkjQt+AL/F1H7x/5Sjn6ZUalPf4eT0z3BRlgzJ5gQprKYC2AjJ5aE9s
5bsUtThnZf7JhHOJ53I5eooTA86utQu0eDvip/NrLLyAL/yV1oRO3QxBBEh4H4cQ
0y5EthTp5NuyuONW1n9BHIPCC/jExCXG5QkLOMlirrxX4Uk3Vp2Za3hyf+JIl0r+
ZtlayuVotpA85Ykk9KeipJKOJOQgevKQ4s1J3klzCSBbxP5gwYeoXlfCK0PwMaQt
Y2aMnrZI596Lz0S87FYhanXRJiac9t2nVn+6LtezYj1WOszSBjexO+z1O3YNu8xA
UnHvlcg4i44otnt9BlOacoShUxXlvA9qD8qM5vV7hUobg89aWzkUxTuPd9vJJzdM
TTxiAApYVis4O/neV7crXilILn25lONck9sT/POjVGX76ihdmKc9EvpIXnLmETXL
JAoXwM396cGv2sD2bOM6thnJGjLZGcBKOMKIHpFexO6PDR0HUc8TYb1XIGuFTbbT
aoI2+83DAL/nVPih7jiEahpeGYMpaBtEOugPIe39zfCu2tLzyG3ZN23RQrYXMJC9
80DdXx/fVzm4dLawi3fZ+t3U+3WHM3DWXFLwiyP6CQ5Hotie3VNhYt6vPTCvBNWW
RS6ym+bMW91VS80G/yPWEQj62XQDgwyIH9RqZyBWilYMWt0A58bjjkI5Ih8drWaO
LvQE+tBpqN1useDqEjqqjItd+HbfmF7XWlrye+EuV6V+39wLs/6X7065F47ZlubF
CGUswtAnZs11PkljtDFZNoWISLnnj/L8syvgxTwnZA3kfsZCHRAupu4o0/8WFdlD
Q/7Bo8u3lizZIkRn1mjD+Dj0RbiuZxYSU/DkpDMQNGu8HyUyX1qwgs0dxYQl6HMx
ia7Mk0Y8tJjBcQg6Va9/3NqcnuU+a6+SeZ3QOd/UoHIHW5AsaxOR7yOCvkt3SyX/
Pqi3HDc1HU6ykxRwkxLrd4JumN+apmph9N3zGKnqvpACnHALSH1tCZoI8SK51W/w
z4DJxFEv9Uhs/M7sLFo4chQkRJ1q9+y5Ec4gfXuzIdjQh3deKVTqZjncHNI3FYFv
d3+aErOlGZQ7RU/OTwKXgNO7BT8II4CoboNdppG5bAbfPJb4PTg14lPeydSMSD/A
b5YISOiP7CduOOr7xlVPBygu4VN2w/+rl30yfaLlQyWMH+25RkshZc/k1UK8qo8l
l1+mfB9FHjHPFXny0I4lamTsBe02m6bfHyuvzZGKFoZp4hl8DxURqEp7jcSBu4hA
rnEWcAseIcXo4QiJ5Fsfcu4sqGdtSV+Zqe11yMDeJXFWnz5zVcfMGdI0vTvWeLFu
oJYt9Inz3d/+fqzxKYXzgv7D1hybc+NDCy2hhKHM+FHjVHweKNbOriq6SMoYhZ3I
lNXGbgFfAlj/yRD0wMpMHBwefI0itTFekYc0iCpR3UjthubmPB2z8Vx8MyPy/guJ
za+N0y4tfbqhkCDw36VsNir6gn3aYVKztZVJ7zzXRVEmfDTFtBtFl85G0lIXcrod
TkS4xTu/yn4U42BM0Q0/X9kO58LcKk3c1b1rNxakrQl7j1zojQniVeI/33cKhLOu
GL06n8pqslNuFA12P70ofYJUUCn3y6lc87g8qo9E2YhgiM07hyeTtySwbndWsKmA
KK99rC9pxblElWAjH7ye58oa3RfpD2ufpR7ZkVfjcMc2PXwBzVGg8t3HaCo+PNIH
sBfvx77FJj9BpaVfvdsvSYCgJ8EIkpQmlgs0X2o4kilIqSDhrtkxOEFeTP1Eb54Z
mFxCZrj/ov88rgNdt5NA5hvWnhVvj5qOYmPJBXZoWzCHvUTzdcRuOPaQtN3P4nyY
tTg983vl4rBuaBOYVYOp60a8pbtdBtrHH2DlLciG0I/YyZxldztFhvQ5xyCYP4AH
Z/4XNojJsZ9GdfwtZSKCKwwZX+oZqqsA0rtbXahz3uUZcplUe9br6PfDEVhAfTP+
/PqHXLzzu+2/ZCmzvEoQMmDGZ3gMkL16VOqVyI/+/de0pRiX67X0rx1HlSZxfIi8
Poijwbq5gWNfjUNdZ8HTLxjhZydHkAJcnlUKJm7pNFGX+2CQXfQP+VXOGrrDwnfF
wpNP6C++KxOPG0AVVgzNEwgiUpsdHKHvgu+2zhDZQ4m6jV9Zj0gIGz9836qT3K0G
WMFzm3uZ778y2rjPtfWf3GjAP3DhitvGN3FUTwXPDeg1RQfy1TfgBT9eu4+T9vqm
mRfwF4nAlcrWktLyHayPaPoLlll4L4ggpQlu3A+EHWFbxey0NjAg1dZPyChOOdvd
wovGnBV74kRiW+wTFYJnaBDGseOn9gHf32bqHq3Wq1hDI91BkYaxM4G2V2cut8ze
0BEWmqvLJShmegNeEbccHb3X16yYVe+lMW3ypITeMm1UhCrggXz8Wr/NKiORANhy
5QnUIuft5KwiXZt340sGp+4gGT7WpRBQ3eQ6HE08uUtpmAE55phe2BzIZQVx83by
nFTAW5s/21mrUe/lFjsm+++CXu9NLnumpRPbJrKtbdlI00UK2VJb8lmQvksyKdy1
4beyOWelqnh9QVIDZMVYPU6k0d79aHlKxsufdHygs8BNwnu9quOVuhyq01KvEPN0
vHTAIXU9ff9N9CYgotsWLvxAcg2nkkSbFDITNBpyDuP0Ir9c3RgLfLkyfulfCm28
iyLFMp48rmUoXcYLeGkiZZP3OvEetijCztJy6y7/zNq6a04GeW5SXfNFUkon0jJ7
b7lhp2Kb1sj9529R9u1s30ZFPikJSFAFyMNZLKmsxAqd+YKrmO/IvLqQp23Hga0U
VNFz0ukUItaqsmvVzuGJ1edYK9LO7zLKRQ+3TWyRTzCxa6dyWMnYNcSQn9HAypHi
sfJnbRbYZ9Ai+6LCc1sUoYaXpQmBz9SB0k5xvBXRG/xg9MC6I5Ed6sHo1+eYX91z
j/bH9MZx6OPWiknWhF2fNR31D5ZYnoi48PNmdsTkoq6NIH7E41wCWMzq5D2GO2J9
BPLUxaNgo2cdbefCdCg4hNuzLBEi1+7WitrqitIUZfIzOt7LIfbAA/KoEYCWIfko
rT451oEhva8a5/tl2s/6TtEGZLgas7cp+qQ+Q2co2urjRFAfZr3JsmVk7j6vgcWB
RuQ7K0FfpEf10Vb+bouvvKhcf1ZmXQl18ERtf9sdy+yAplDBewNCTrWjVV29Gq+V
Hkqqg8i6xsW4EpOwqecPb0ItnuyP0WHXuuw3iq7/p+gvIEzPuz6L0hRZWn0eObnt
lsezL2uGXr30+6YuYsmRAakwUqIKLqpgxPcUliOHXotOsZhxQRzWdfZOl5dKLru+
c22u9OXtFlu+SZ0m5SR6Mx3sl9m6Sbb1b24A19FTcadOE32FOSc513nkMUyHUHux
/hNTg4inf8J1r+z/X5jQayhSVWIx6z0zQFS+uQxBNaF02oatkY0wzCFbH3zJ586r
I5W5L/qELktEAyBrrBCWFeRaGYpk3+jFQa17yTuqPy8WJAkcPIejgBQ36A4AHukY
oHTspuaQDs731dPJNTXZKII3vUIcv9bXIsWreAenkZWCgO1iOllYUYqOr/AaEzqd
Y2IxH40yjerIhmQA+tUEfjK6q5N5UwQMX02/zwAoJzW7spRkMZObuHyR+DJ+vjRp
W2h4mGA28aU0AsNX/fqKMtsDdciLRpdVYnt2yhx07n5IP/SI4c8HUJajOj/AlEWX
0m6+VHHc71Orz2o5GEhs9xwc43CeYrY2fP/2svBz4urXbJuAuK98jae/+NK7SnYW
N18AT7b29msX0o2M6ZfdcmGjPZ+mD4g/2jDy8I1g0hz80cljq3BswrSWSe6Wi5iS
hEQPXSrNIVjHtB679dxPHiUkmEm54u/yFgS0SuN1lbNyeQNpv8mTj5WQAJ5UXfGR
4VDzXPWvBUlvEbCCd8SroOL//3TsnS47ka1Y6aNTT0AjudxL+2Q800SUdic26MaQ
IHYMetyQAfHCHUJHq0tFnfrRAqDS8r7L2X9L9UP+76bOdnrLfTObVNp8sBeu0PDM
MGtZQycJS3rvHXcKU6tvBF4QnG+C/b5uNmuxnrrHKdk5WwhuDZbKFmPzz2Gl6nVD
gL0eXK+VD1CGyU1fZS+PRW79V8tHSpkDIkxxx66M+ThFG+aiCvo+iOcxXyHuh6sT
stnDsI0favYl+DKaGMxCaOxgGllvyono8BVpb94HxzIF1ANYcQEjtT3EfKVMcrmj
3M6LJmg+rOkbgtV6Wx0PYqZfG7fYLzfeszRd3QBk0WBX03Cl6+xUO8Lw66FioID8
tm8s7igfm/WgQb6hZp6XKToEQ/u9i0NIjuBtWu9Cq8bc1Q8U/QMOAwt8y/TZhQQS
Kv2Ka7Exzrw4kGER/6OWn6NmUmkDSZtY5djOt9XNXHzGODUsHt6JWbo0FgBmdZbF
2ZmGcEWz1w9s/ensOVOUszWOhNvRFTjRXQihDZZyQUUfxtfA+P3GnlStxM277huR
MLzLJHSdd1uY5hK8ISz0jxWmp3KLV/oNHr7z321oxYmccoOWgp+jNJUkvxrqO3Ir
m4b9hXqD+rFcGy7nkRJtGDUNEcuE+HibjStZx3w6wzh+Hpe7F7cBa+454TSZlDRa
JoS4QcLPfHp+x/E+k864z2LxcDVnUqnTVOnBURbS2lblhqrDcQJ1mXny15QZFzud
qYj6UKipxRJHezDQ3A2Wdx+p/BT2DCqtkMEUpgu2rInwpuZc/biiLPMWpdA6z6Pc
MPtRo/sCtr6jxoGWgDdD33AqFtXat4XHQgj2YctncH43KSz6RcKt7DYeOI0E04oZ
cguNJNY9I4RSDxPaEZmbgzkPBWLqbZp87dHvPPaopzsgJGUm3lpNC1sS4XCCqY1G
Fb8nK5ue3ORypewj9mzzsntw14eL8uKwJwnGj9lmHu1gqF3fv1fY1GDDA6NlqDLD
9Ybj7yiQYiLijBXCNFG/HrnimpMVSLh1oRrJJb8QRYiGA3uCud1J1qhkcLaMxbBV
d6Bw3n1ZvKerhhxZqYJk7dcKqSfqPy6Qxp97MOqEjs9c9HcNCk9cty28eY2PpPo3
9g/imvwwJUBR0zVwq8XiRRAJaWSh4melgmn8m8trZy92Lr6k9D3NkWKTW+rcd4pJ
WCxEMOI1HdXp13gkSjcMj9kMedxEEg0s5By29uuNHZGbcn9EeOGb4GDvdZHO/wfC
CZ+CyI1z6AgeNwdTmlzRlRrResnh9KV1s8P0xslPFd8mX4RXOIvpXnj3lRTkQQ31
WrFRLJHkJpwhcGHuKFiDC0qkiQU2FG6myQUg0RduT9oGFkEPUK8ktnYSlnAPSPty
TQJkIBfPPMLHE2e43o+ZarTI2dfGDC8nJnBYrBh92RULLVx8knSgECjEZQlvrGWK
p7ULnWVVAMd9Kmy5Y8JU3FDmx8QAirkqU/KTIAbD+l6vAVKCQ2FCA0zfvpBczRWV
l5nsprcmvRuADeMiUmh/zN0BqDamViCvs6TVQp1Lmor4ccXzf4OLlMv/Dmcp/FrG
hLRUAdPqw8eJp/3PNcwKM0Aeb0pQpOQDZg9XVYAEZJq0AlfyR/syazbrrCSHLd8c
kgPELMvIGTcPkZUGtBnNqH02a2uh4wNU1Wky0k0bnuPBson6bXKCdax0tE9EGo2e
PEEtrcFW6rsi031a5kTwMKuN/Q8QimOTnYX9h2QlQS3nwo/dvQmVFe3UTw0P3MkE
doL9AmaLuQUoR9bfQUxDOw5gfEloOKueFgoOO4uw7KMq6wL6SEh+O1/4ATTFmvSs
vb+aJvCURTTIbtDjrLb0VJDKv3yWCoVMYlZNPgdYUXjSku2w/Dfi5lf1VpaL127R
zNm76Ey7eAau7bAgi31fryouXqjLh4ZI7PcP6dsVWc881PYE1PpXccLSnWjNdYY9
Lul3iW8C3jkSimiBWNDVxjyW9rL5ihh1SUREANjbrT4fkPt8TX0p9tOgMQCbWZWq
14U9wiTL9a/RBQMZ920HM8/z/qlT8hS1ILfYNN+3m33de7aAIQBvLhVPsVqTGaL6
dmlb0O3HVz5ilSuQIKJBamIv4zs5Vo5jfgB5zx5HLF72+hyBHUBr/mo5qtWHMsdf
NztnkyP6Rj83v5/yelXHx1T9jMWxuV0STu9ok0xPtLEri5rMrO+hVBBSP/4wXQzG
ug9Y3iyIhU9++YWletx0AkJHZjlljhqtPt+pTFHUye9Hd8uE06NU5bpwtncqAZ8u
jjh9q+ZGGFTwuV0coadd11I0Xo1Sj4lVuIm/3JqWMYTLHKwDXQI9TpxF71bJcc7h
/ua2djBSao5rVnkhtKWWhWXhSnL5eRv9ug5nan1CFxVZL9/KrbZh3yvKXILoumlA
fF/OqoI+q7nBgfVfP21UKCMtxnfUizJlj2Dt1/kocGwzJ58aeFjmHVgr5fjb2aqQ
qGtjt6MlifdCSGm2Zqiiadcd531Z08RCOy7/Mfh+j4/2Idd1GMNfpYdH+8bXAsHz
5C10o+qsSvVyg3VPW0rfYr7XREr4G01Kh5TzQ8Yf8QIr8GynofHyiQlA2zap/ZU3
8l9OqbGIryaCbe80Qp/mjjRt57XNx6LkHToZo+UGWvYHwvkhk+0IzbhDZ30RGXhR
NLkTu9MKxPnJrtwDDL0wVE+T8CakmaCnXQL9NYIr1mA0dKiNuIqNx429yX+dELGE
98C/NS84D9AwXImgaE3oDIjbBhrX5ynFXfKR45DgbZM2dNDM7sl2v30wnp5LX2uL
pS1no3nGzQO9WwiVMa37qZntR7iMSPOVGPMewVIQqTIXgVV+eT2OtXXRgbpZlBuK
HBWFeGrggfR8B4JuQGLpANiMIYzhgGCnxirN+0TORX15LJsfGnesRMhFVTLKJWv6
HQdO7z6WzOyf1DUBmyjcE4MDrtA9O72TzuQusunUe8dZ+Ii4C5HOp0LBrsEi0uXO
bnZ55Pja4WCSigsE1CzJL8KjBQ5shjg85KVNRzZTCLrUvQAzt4b/it4IRwCnxz5v
HiU0aNP1rWQKw3O/dFBg6NGKMKhtRVNExlTEt648phJUMoFLGlkclcsop8p4GMnb
NugI1V9rQrdPRNKPObf9Uj7kyeMxfvXQxJFxmKsh2vmVkUi6NXh4bTCGshQKeliC
t7vDNonavSULEao10PixljKRXsdKJ8wnx1/vnk2bVOh0340NE/LX9o9t+luk81lt
GaCmfKTdnhOs9oiaSO8dlsdy0sIm4hkSiXjbPwOF6OO5V/c5nBfet7tmi4A5F8TH
K8NhMDHRVuSuWggG8cFcyZCUq/kCstwU2Dv+1lbVOQ95hRrgMsWGfHcg585cBIFh
A02KWPnUnv0Q+Xkytf/3iGc1M5FQzt8YqgjYDkkErgEAd9E/jva5VZfhyKPLDJyN
N3ARhKBl7qzNWpKpBHrtjIM0nmf360hEKP4o5uB6l+0tEK1Wu4yxg/hZoZ2hYsvG
ICun5ht3kKIeyLeVS4KKJpOdsSdXnVClZss1Uy/zFke08jOMWQkQqOYdfcSRNm1j
lF63ClTboDhTHZZxCVNHo/UPZzVdw7a3TlRamYB9nfIuB88P7Q90Q1VtOIXTzT4t
jH78m1HGkSM8Je7znzijryI6jzWmHwOgvzhK9ZvAlYO9fz+2yZrN39tiSn7LVxmY
J8HjaUSXHvNTN3mPJsF+Nv28JfGUf3FdMS5v5WD1AuzaJYiN5B8IWY2LStp0GChV
Np1MW6TJY975ghM3WsX196X7ZZZFGGxgYcPXaKG9lDzReqlK2k40PLTqHlVI6DZ1
EwRgUbLgTtzcSwAc90wrgGF7q3cn+wvpUg6h21ztlMKsc2pzyR3geRskJlDUCfVY
HNph6iVErw0UiZZkrCIihKqfFYR2g0G1hPq4Ta8TnPRAMTazPLSmg8yTs4SoOsJX
2jliAhTDDcSuLNggP6V/V0RVgTvnsdJlvuRAZn1zwQXGXku+MzZdg/5m84OJeYz4
7gMuQI+qFntBVgT9lnVKWAm80/s3wBRebbLHXTesbWUYlYlOs7kfuFFp0/whYY28
KD7fWqDc4xF/AmcXTBoG/YU5GN7b0JwKcigg7fm0llCNYeEJF/DjyE+XdLmNAKNa
yuYw16geHW9iNi5ah2Fqyn6o9VSjvbIdseA9/IcbZ1QP5fHLhkthJrSoJA4ZFDPC
hkONpuFbaF1oii5vbMlBPTn9ZM9KVcskDMYjwG3b6rsfZXK5FTakhWvQLuBJquyi
jjzR3hA6Z/ASbZBO3p07neDzUcz8rCZOXMx6uLpvjP51gXDUhWTC4cMM9rvB1ESv
PQ9M3ubZtKHFtzstmMZ/K6jgKLKE6ISx8SrxBj9Ldkdx+b+0vS37hUaXhlcy8yn7
BdzC3CAM4AlL4zhFoSy85IUkZly1/t70/+ghh8AbO8g4vrgiGVx1pYGGFJSQU0E7
JohnL0guFm7lOn8bk26iFCJuirPvnEHlqzQnR6GLOe3BlxEGXV/mXLTqeDA9CFyd
8qzoPR819UE/qfZWXQkbi9kEd9mSoH6Yy4d5lcGqjPFGqqKuuGtK700vXFbWkaLz
MrTHt6sZeigY7QyKCOaTJmo8KkeNJArl1w0cVgi2HyFwcQqOVVkasIgbB0Pm6Q3i
vFStXGTYqPGyEN89eixYzR7y1uH24vQipWkMuSdNVaUyZ+ZtJMgML0iNyhPcm0TB
qWfQ2s2EFHDvIvC7qXc17m3Nq660dga3EzdQiYgfqifU3yx+i1Y0782VR03pA9sZ
AJQjgcKv4iheUvFbyRokzOEWqiYXe/DnMco3YOswl7TclPjxrG+RnRoGyprqR+M3
8Jq2jfjqwng9eAUt3F09e+zyRugV17h/w89Jrr/HCOPHqFs85LZIUiCk9kso5o+O
v7zFY3Wd0zAdbvS/aGiWkEG+i1k9bSBNQlRo/Zd5MGlq9gw5PMSKzAjgoMv5EvM3
fzHlm4cvAaDTTwPyRAZz25g1prJ2H1x5+/Jt+Yr3regO0DwA30/EOW1yAhgtvrPq
NBQSWjV4TnScN5b45ssvSrisGB1Nv4A7bscMM67meIVJEAlATAccSOiYgUhFLMic
dOghST39vjc4R/CQYDfmP4y4GP+oKc6mb9x/qwidndEHRbUlCHmb/H5ZvL3jfW4D
AhuNBMPhsYuk2K6B+kkbExPDqYrMV72eXDBUMyHRcD2XZhsAjp+8HDt6/lkNablx
v+73sVQ63ZFwoZMF2lcu/G+hgS0knubhLak0xWpZSDKxjZaiQWx8g06YFH2bEVVT
B8eUTHbdYBR2eqXbF85QASDLAc2e9yf6Zsk78eyQK+lOCUowhhYiYSHL8ogvGnba
c3FauKSOgs/EC4d2EAyXLD2N8XZpsT+LDAy1Py/x9REfKyeavS6MDjcUpuOu+NsF
2olSqg8zbYNwrhok5vygfWcT5JVV4yqJhiy7s3rerFQNbDTXnY76aG3yQ5UAolUB
pZ0n2tuNP18GSQ6tn1w9p5j/7Os2k/RtL2v9J7XwxT9Lait67I9/gJzAVEe7H/t/
1EnfQIRib/HNpygDMnhLlrnEgv0uhEs9fLGZaz5ISlHWAB6+PClYFi5HndaEjZ1z
slUK1gHXaGYejI4rU39JinGaFwKRJF7ddJRqB9m6+TVNeqaGBxnNEyLSSryjtxFE
eUcDN7pdACSkyH4nRgMMa4dD+r7DjNQ1mWvSeJJ9sFwf1qTt5b9Jhq5u3DDB2m8E
jh9MSmjamhv1sEc0XTep+bBc7t+iUum5dGM/wdy11yNjbv0EK3lOkC2j9rOk45vE
/bCHO9daK739anha6xo0MjzKNja4R1RCvIqW9aEgWz8BzZETBWxAv9BLbvzH1Nl9
t9LdrDumi4w6B0c7Ito1lZsd++xPTEllvsTe2AJOLhSJn/+fngyhukxR23ZC7UBQ
bFLrE/hJUDYvAI8JZi/5OnZPjWNN75aEx0N0FwwzcutH3aE+dWRMU9a/axY4+dlk
/nfz12sXzDlCzfASL7axJ73KnBIoZ3z0aFIvJaQ0z7aX4+kuRSIg72NrtfiDN5PO
2+tlAIxxh2JbGu0H2TU9I7cZ3XSMM4jQsLv/AhidHj954ymt4TvDCo3xtbAFgmIE
UlxaX1pTLQGjHxMwWRMMEXKqGbzi7VZhUZS2sZAgX2k/+VjAt1M5FcbUy4TMPgvN
DgBqvJN6OUmgnRYmxOYXtSWYd8f1Dopaq0CQL5ZlSyPXTO2zI6LyoVorQCUaT9eb
BkZkKMMWaNGQlceGnzpfNi1LNuRwfId2SoYAva3hMJojpLc9Ov6Mz310mYzsHwtp
b013WbRnSwxUi0nZRJHvc7a0jGjyHuSnadCIQE4bFH6+IkOyAf/7hnd142t6f2db
df2VfKKyI9v+BzJUn+pgARXlcEHYZhwfW8zMy7GRNjLtbZ/QEEFv6KVSPo37JCVH
bcYLPjCL3Q5zrA3NKVIPr0a9vPA1lIswQVy3jquyQTBaIQMw7pQTEvwfCalWSJW+
KeDrLMGDgrd/C20HF9zZZOi3Y5ajtEmICJETPiFRh0U6y4m82f9rTJzukr6/Ssou
sWsAof9/G+Yf0w8ACBjPNXIMPnDir+hGJS8Bd3fgkFos7Aq3SJWcpZ2HHFDFOBXR
qAZgpdnnTYNYlTfTtg4AdwgJRbMwzH9KWaf1XE3ZU+FkpZ5++DYUgFAQ2qT4tOxs
8q7+JhsoCCllVCuvdNaviZtoypCl+m+w0jAYN6e6BaREmXt0wo5zmFF0nw2ZOMqQ
op2Hd7q3SueF+ndWHgvdqnXzt59tSR/85WZxapYItO2a1671K3KygatFaRr+gbpx
UHEfqoUKKEloq8pcHo9auLC3TWgKvJyq18hFzNaRh3ZKwCOcFhVmwNBBFGbiljpO
AmyskUcSWdft2q1y1CQE+BTGNGB/RiSdhkJk7sgw8d3pQEKmqIO+RkxWDSLSG/Zu
hsxWWyZBDdEsCvTBEpZdbnHyDrWTkGMXpOG4jGNz2OFJjwGiGQfAAdh2IMO20YNj
y+AMqBdXW8eMYLIBtzZ7aa1urXpHv/HTB7r709CGP4c/PX6EFRiNnt50kKWV3juU
DYMTNY1oFRDv7R8nWWY89EVSVHPlPfBU1l9Lv1c8S/EykAVno2rly6vc+ifHUxRG
4FeXLIm1hYaUjyEN16maV8V/TkS/Aj9NfmVXHx4ZyJdvBVm4R4B+rwlc2QeQk5GU
7zQZGpC/MkNpJEIgMvIZgi0/1fhD9PCyP7pSUsnqx6PZ7GSFUBb4mYxtMkoxDyeV
XQEEGphpAeVpF2vBQBN2OARsVqDd9UqoXGatl6C+5DZ6DOKY4IEo+yaSjijeIrSA
dBKMQl961omkfMrZhsbGsNWFiNykJvxVxtY23+Sv9NxULHItXaaEZa9O68EhTgHR
BqKRZzHAwS4HTwBGs/niIW34ecYEOSVBccagShvC22p2CHxW0Ey/IIo4Avs9cV2G
zsP3YpS+ZLXkJILXB1CnDhrAZmO7JXCrq99p+DH/DmjlomEAvoBsNfvob8oC/lIE
LlefaopbGRmz7jGOBlWZqxNyBoaRQuWR8CWCgAT8punf+dWMvqMpHm240WKZckEL
kIbPTN9oGi0oAEPrPubnkaIE08piGS8H2W+ekWvIcQ6uCj2ZzTnW7wv84MzWcr/8
geBjb8HPTMPX/JLwdJOWB363UGeGTuhErZbga1Ma0HkO4D8JkG56h53YqeM9yxOu
D9HvuAGgRzVqAqHiMwrGm7n/K+CaUZJmxckkJ8oUBYFlHETjvXxvg93+1Ciyqw69
b+R0D7eRln9T7UX6JBzxIZNMnpcCypdkXlJkcNJ1yVzydMEETTIFi++b5D2vjgtY
MrXDz50P2psth6xtkmHCwSO7yfG1DWhdqKOH9JKSdp2MHg2gp5oSQeYFqvzmgP1o
x09seggIQ8uGI8+9qj8R9+0XFzmxETXec+gp21HUKcya+umfEpsJMNdY6iLyCOmQ
M2uGIoqxb+8teW3E0nYalE1+oKCbys/zCH9i481XPH3qZDB3QThDlLaJD4cAdYXP
8DUmTaI2/xso0gCg2yZup96ztetyZD3K9Cz01NdlN8sGlQEc8NtQIQY0jL/LPxr0
4OmhOXLDAaO+NL6I8LP2OdBVNbuFFVa8E23zdKc+T6XzthucwecLrYWtZYpaCeEt
aBqCJwT7rzEkflS78NvCd48y5s7lpAYIGoPsHBwqwy29+sQkxfBqiGhMFs4L5U3g
UakM+npd16T+Mdk7+7cO0mStv4krKr7xGqrcagszDsoKD9HuMtpm2wlzGxQWIo8/
Q+k/kYc1ckDhxLx2nPxE9u3nz+voqF4RA+YrzPjEYjshgYVXFWK7akymEq6XlXk/
CHRFBZBdkGowndjY7al83GZxNp6Y4mjG1PQXh2GaEhHCN0Xnf7W04TJ7rTU6s6kC
kID0GPMEYMa4HK/TLYSsUfQD4zMRK+yMiZ9BZ1MGMuNqeRwXVChaC3HoHicXdJFU
DBcghwpkCAftL1Pcsuf8VtD0Bx6WXEBPHQ2Y+dU3H4GA1NybXx52Ax5VQnXLjSIr
FQua+0efAp9CPoVKwajNWSRlInIot4UncRPemErPkJ1MIApVJYZvwGbAZEplwehk
C7rxkCyHeqIX11SUTL/MhV93gPUjlw8uC2BLiG93Kq7byixIWactX5vZvUZc1h3e
V/k+JydkX33ybFBPWGbXhUlMvWop80OzJyeJOsYIxC5cbCePzYOHTDakZY9tFvyF
5AYcEgy2WNwLwdFYVTw3TyIaeoxxcyOxIv+6Qpp33poB0gLvVnf06DCt5TbqYVuU
ottv3uB/BsLHuaO4Btw/GyHaY+JtG7TVO7PhXxy8+ZZnzS38ug1LRMnLtjWopJ3z
d3r+soDkla6cqE/KmwxUH3Hvex1G8gLji8sJ7Ejp/Cx284ks1WY4wY6JH4b36NK/
S8A4e69DCRac9yF8plnJ1zlaSYrDKjKcXEnX/oK4dSYdtdmvG+0BODckwCmyYhea
oWmSPTiqljFTaUbCvWyiF74yPC7muv/U8joIX019lBRol46xoaWOTBLIAeFoxgTC
l15VaDhddLc/J3TY9N0jv+UZEv6GswB8uXkfLbPwJtYz9E7imeOfQ2tycuw7392t
DwGqu5BfWrOUhR84DUMbX6gYjb08/1liDfISmBHOkgEE4ltNUlnLUgM/Ylbgfni7
+JlAyxfDGnMeFDUrJtSJnJV54BYXk8OiT9OPrxvcLQ64rMqITR9OEUZto4gwJhNv
pEWBGd2FKBrMK11DpRlOq47dPqJtDFyrTZ0jZLiCzCavsebmuWdEyhYGmn4VO6Vz
jYAGR+MSp3uoMJP61MVlecOAKDD32wWMTlt8vbbRkLz+U0Q4gSohsp6nbcaHWDSt
9FhFk5oSgRjCuHQVPJIvRBUZafIU+eFZ2/Ku6dYJfKdf1tg6IDooeNEJQFPD3FJu
YAT08rB6ORE8/jCE/zdv5xyRrRvnhksYvmnKp755u0ivaB5GcDTR9pvv+hkg2/WE
vjMzO2q9Ae0sH8u/kC2vFpnu/eGy1Nk1IsLCoI9QY7GP+00GsYF5Qj7dmMoanQ85
5Kd/dl0oWXAkvMjTocGF11amVyMbcG8mWPFdaiWWmjJjC2lHxg56s2654HOHCBQy
DqevJVUfK/CImWpEd16GK0/kNetNRF8opObxYlfetXRO09IGgqtPLgGIrLi2eEX5
MMOwSOWWAoXQ0H1En3wEbuAmLcJSuQL9E/kxjGA0PtGASiN/fpA5WorQ+SNAjtnx
bF81n1wzo1DlKkY+m5h/sQyYoCKwEVJUoTbXHsx/NVKtqdXhY6aKCu8WciQ/OMkH
xlPyqMk8fk18actX5Rlym348SQqV17XcH//zH68cOawndIj7Uh4V7UTfRWxYGygW
ShM/LvfLGBoihjfDeLcDn0DU+ke8RaxAZrpSFsb5RJFPZSWfM+2FZF7gXaOIRiQ1
ta+g06RO9VMNJiHL7bEY+pYmhZJ0W4dAUjgj8jFILGeWSyNMzWhg1dvfs5V6P4xn
A/1n63PoCDF2IlqmyQbn84CMmqBTNv7W7o28ejx7+L/oyhIGspVaLvWwuOpwAaCQ
4KHY0nNQ9236YdnOKFLsg4iKFlNAIEwh9eN+kRlOzdqoPNw2sEc1++9UUB4MXF81
O/ZWVUrvkzyGKIvewyhDAI36f08wqY9AQq5J16bVXEceT3lwwcKgjP4ncBT2vzjH
RC8FOR0IN17lVhtVOFFz5kYGz2Dc8SeEJi6CvnU8EQ1b36YvZWcuQ+fY3BAO5pGb
V2b1hW+/rgsxdZU/Lr3HwWCF/UX+fkF2HzyTBV8frRa3Iv2Ru533H0b+RGl/bTBR
Fd3s6Sn0Hktz9ONvNKcSX1a0XS6sBvIt5sKl8dPfNg+/xb3yWgCd/rvk6t8EFbFf
9UiZ97EbO5tRHtcbRLqZN+wSC/PSKT6vOAlzpwwJhdtnEJe939PNWVbB47Dwv3m+
xktms8mYuet+wqXoAjSVGjGONdaEARPEVKaw3NS5qJTudTPVDsQmfj5tf1IAPTSD
yjsuhpSRfI+KIM1U46zHRummenZDyb7XGbQVcsPI8cYAdNq/OmamuELEiODrE9nv
m/zS9kW8cioLIEf3rbj9stq20W/55s3V5e9Tuj5OzrsYkQtdOHYff3EP2cb8jN3A
TUepcnFuDsz/Z8xTz5HO3tP3txhREe7sJAAXGHYj8M6bIEbXn5QayGAFuJzzyUBL
yCfKPaf0Ux1mUXE+3qzSBaclz/FEDgZWrfiKi9x6p43wFx3UigDIaNFLpN8C7l6v
B9pycoBMcGaGd2vfmANZ7/hp1JzaoEEr7TmYlbI0C0j+zTR13ayfoVL15cREvhmm
en1XVciz6gTQPYDXB5kYJpXqK1gfYc9FBZJ+Ukl2UTSNDwA5uWxbQib7g5ul1IF5
u7PCbsJKXlgptrMV2eFvQSzAdQO5BxyeMiuHLZGQuIQRe5sqOU9vRSsFq73Tyejp
2vqqXyLTSoHbxZTWqZzzZJZ5WIFj4pirxvpT1JNqq1k+Mwq9etbsEmGgM7Q5Ruww
px4rLV9Fak5yQYgIV73uyxg69SsuwZ/Qq1s2uBEjhJSL41EjcsYLro7KHeZBz9xt
NSCXXitqVH929Y3eDldl9tuXbG9Eq4M/sVM/h8XY0cH7SP/4WK7ZDqmyKpMaBqFK
vuNHkJWrxbZLzRafzP8RNKLyXR20fe4olw2jKSjWTaYS9g+oW1Wb9ZBJUKZdd3vR
Q8eiED1pxSQCNn4fvAwY8MKuBiKXD3loTV4evZSvi/0zzy/ePFJFsS+JM3AdPdGy
xz+Utgby9uwDM6Sa8jSu0xNg6QGp4MkGhunEbK4F2vhSsqeJmOAZyO5su6eqiZiM
S8IYT44kAR44SZMhLiNaPmkZzvvJOpus5VsJ26Y5kxHU/hz9jZFCgUoWjd6tFlR1
jx+k21I68gNWf1249pIspQpcqZBzMKYdpUdkO/+L5NKFm3Ntg2UeBwhJlnYI/0l6
4wsEhhivKmFn6psFnSnwqyEURMB/xLlcpmZdvm2J3NCex1a2oCgemtfb3Q/PtP44
sRIsbjpHfgOlmx+ImWa/0TaVSm3xK+HeN8uJTZKQopCTimgfBejpZjBwe/eSqfly
e0gGQFgkpPr800I5Pearii2o9CkSZtE+qSG4n6YkQ6xQXiclQhZy3NA5hpTJDo7c
kzegYlnaCuAFre7pymv1AIemo7yoWcvXGWnDanfhQEtG/XCmqbSmRkuyOWqqubFd
dVlQZEYZDnkKCwadaAfqocJja2kWjcCSvJ4t3xL6yJogAOfuRE1lEyj5VBVcOR54
E6FKONuw4mATH4uH4DxwgIB4qEjV9IrImhg85aR6bRs/lu1w3wUm9MA/SIvLdOtm
r5UpUjyXA86M8W9mwpr3uT8Y/HcfD4QpzdN1NeV3WRsOSZ+1q4CYLiYrTQXk1Ovv
+wY/94/6SA05DU1T0kSiVbA/LsIeN6wWMjo9HwTxaYaR5CkrHzr0d7Kl2jNynReh
1O7vR6P6ULLGaXphvxeJhyIrSgNo9FqUWmVYPsi3Nk7VkH16ctrhgQKgX/wKCK3+
7MnYoQFP3l9Zx6Gpgd40fRsZtVoMIliFfLpUoWD8Dpq7YRt9u+Sk9CTTSqRvv6Sj
DyBFQ5dkk4WehxLgLz5iqd0Y3pP7y4NqE+V84y3SkHIX2ingRp5jxKUSFzuGVxRR
RkaOYtsiy+/axYvURQCvjpM2xFFBNwfV6yILFkFlFbg9hqdYTazvBl7OlNcjFey5
0S6gLloPlFKFOKcMZGDcKbwsgGqKv30v3A9iFvrpj5th1WPgSzBPZyO/n0B3Lgc0
1US8Jqrgqjjkha2h8Lb4WrKMOxNpKgPlutPgbzW6fEPG0CoLEQS2r+CVmn+pcvfu
bkCw1LS7L2OQhLzC1A6cX6ToUHR9OeeRv9JamkS6jvvku6K2x6tNfb3OcgTqIM5m
E7ayJ6QoZF5jylJr5INNYyIuj6Dc8kahMILiTFFPCt7bpqrQStsxXXF3ROr1jjPT
1XCsmIaH2mp1QHTG9occu8LBIf++z85U7Rc4wbVpuyP/cOCB+1/RECgLSHoVMMIl
wxgF8/Wi0yNbOIMoL1l+sIxAVKyNB3qkdpPlxzWIBD7NCc7Ts8hR0BOrQHArHwGT
wiqMfyS7tfGG9dk+UCr8616a4qrC5C3ZcS2UaqjXGlwZ6Zg3vNOwWdVDBekhJgOc
dbOHviOIfpYWs7HqPNWAtodclSRguIetJqISz6hYB18gWYQD/ewS+kX982IoujL+
vHxmeR6U/GbSrlw8EurImFyCdJGJj9tMS3RQeAvp1PrGPHOJo48TNNiTsTdrhMEz
7BsNZ7RGJjk74j83mjfcf1TiOFo8QmGPABNy/7z7+HMfYjZSwIYeLjtE39lp0yMR
JwByUJE33HiEr64J1K/WpAc2W9L5dS+O0sBEtbv7FE3ZVhtgpFCXtVXABfbz1x7m
nQaO1XaOkVlNbWgMY13a8pLt5Eapnfz6kkaQ4WarKlm+hSfsXDKgJK76Y7kQgqal
yBZabSbrRLkPEyYLeKDrtu+eb2+NmCOQ+v8LB/0NRPq+Ifarngvq/lwlUE9ll9Ql
bcGT958tBiOPCnA2Gg4QOUGhIRh1BpJWi4/pbys1GhK/P5TMqKMo2m3NloEl2dui
nLL1D0AlABThx6HAkkFd7CBYLsUnsBif87Gnq/jtZYWUW0WgHauA/08rVHExDxHm
xcj5ddku4owGzMjMoR6PoKvuU0oaPG5+ONutuGuCrKTyHk/Z20TE00eDN57CkdgU
XRfBc/3T0tS270AohuSINAGg08V5oR6Tb4pVYXhbW6cLgxrl+333NZjIpOSajOvR
7woA4hteasSq8luWSm1bv+DPmslcr71con4SyfMjABZ3zxI3sGfdZWOsYjszkdEz
uLUz7IncOYu4+DxA7IphHgHcG+ksTkR/6tJ3Jrhp4CGKxmAxCbkNQNSjhNZuZXr5
1jGvwxtg0ZmyqcIRlghe+t34sb+vT0AOrd/SonQYv1pX+16cKyQVCsox/4zA5NR8
S1f7HB4vV8B5xScNGbPvv+JSPFOlLL1YK5QgrM/PwgDTNgL5Fd9Wuai2S2EA7d2L
ZCOdVwL6HLHg94EDpxt9u/XFoBSdx5VBDnoX8hLLjmMshFbDR6cXslO0hjJ7zLML
buFB7UzH10NxX+mD2b/kHcwhIVYVy5bEZfcPXKRil4fUhrDZT0QmAgtjWi8tEtX4
zR06I9Rd0qSIx1BIx+xRIYUfaLPrA3WnKoZJ3Kh6b1sPz10916ZthV466FHO6f2+
c9XNc5G7yA90sPkXAoD/qBg5B45V1Y36yqXSP0rdWr2BuJaq9e2pFA51HtDsuRQd
ul1rMOz1RnFls+ztHKAE1NqjKB+0dRwZMpe0VthnD2luv+1eYcyB2vvit2mgfEnu
LSbdSVzbQrxVgCz+cdo8lQKJbPXdODScghbXoAneCPrFktcAaqFj+LwzyUGs5fal
ldB+gYVXl3bx0AQW+6vNKvRXkl7Zp7Lfp5OEUZSUju4dXoBGxPqA5Qn3C9ZtsfOQ
LbDprdYnCGOr0RRrEJCodzrGpJc6Q0UhHo4yui5I5eKPWf8g7ISNycpwHc5h1CWf
2KKBW0rlbRWgbQw+Ak62pfkrx7BciiDY92PmmZFw6x5bUWgpKI2b03Gn4YG7H4um
lxGLf3Wj+ksxqrGI49wbTfcSTadUNToOFv6VqpjQdra87C+wSgemGjil41jo9kGx
kWrvbHCwpt46liYbzmPuiuOWp3vsLqjHWAXzcv3pPzwdXZsLyc8QzriWLUMYFZ8o
mzwMBPwIQeU2E7m7Zs+tyPdIcp2yPsHRpFEngKA1/UrOvZoF3/rtTNpzOC5uXPVU
qw6BisxIqtoPkrxcDksKJXw+iiISTAen8KuBh04UOc51dN86ELOQz2OV+SjnQ5N7
zEl4ji2qlnMnr0W6joI6FyVw6mZkliqyYWvSDbfQk0oMyoneoimdaFRLQKBLqsO3
RWhhK4TuIdLXr2HC9U7NbaOTLzuZrc0nDNB1UUR1BOuWNmYH4Lu4VQyQKWKREGpC
AUSrDqtK0R7QbbyteltKmgSehxnCKa5BQbaoENTu5xVjjmHzSQjyb5I7H4zxTbcE
Mkbjvg5eagwZ9ZLHqo/zjgJkpomowQR/S2SGCWWNsLBt/Z7JuwcFtoW0Kt2ENQIi
4fauMZR0BbXRJMR9dqtM3aT8fAl111EHfCvh7kKKcmgEiljfsBrItotZE4d2LTdU
hCbdpTttX6C25tWzGR46A/BuQ3MgPm6psj9+QaMQNqult596kIy6XCUiGJMXIuMu
9P3ho4xyfcbn8UihdZDtGqblaDKGnYmZ6uJDQxYDggzwfJmBjPHZ/Cuk/HKkcwYs
Gh9e0/3WZpRBY6MIdPxdT55TpNpivso6YcJRnkKFDgqTI0hOK28KXjPnsI1FzCd4
FqK8yo2FGQAbYeCt56SwLIZBBHVJDnkD8Gpc+Qes1yIBUGdyFfJlBb7Wbz97+YMm
K44IX0HIT8akz0TyYHfmgNsa895dc8NNWPYAXrko2vnr5Kv8Wb/4znBtZvhEE8Ak
sl8iX+t2enm7AVp66IOkfHM8CbfwJkyf0WDeRBbpwQwyGv4Jm0hjUQRhW83tgNYh
WOiPXcTP3/7DyUHL2m6or9LKIo0bmrp2XxUEjxEBI9qLx7Ah0T8XWcS+kr42tQjb
ysLIm+4JE9hfy8e+pGzVEaQKmSI3MvonK0lFZdob4PHnmBxZj8dJ8VvDbTz1jze/
aDGIn1QpNwifCHjoo/dUQGiqaeTf+qBPvGp8s5I/GkzCRcECyBYkVr7mSlrwzqf8
hoCtJFZK5ZKSY6FF49B4aW8FgQretBrB9CXZobHhsENiamzpNosUMW/YS5w3X0rR
pfb5lH/T/EO5PdLw+BpTwuiy82xiSbj8PxyKhuEi4xPT7CrPA0mVq2cKhq1wiyBm
KrE2affO+R/j1cUwmsq6JSzGcuauHdvUaTBuLfuS++S3w3fgxg0pcivW8selyVpu
LV3a4rsDtke9a5FSSNCY2150VLhK5ndGAyxkA9gexA09ZdSzxeduJQzLBXQnOTjU
3TwiTqWHhqq304T8aM6nm39jcASd41sbZgGUhcgrxCkYHESAtup0rpL11mpBu6rh
y325lvXDYdVFc1QQGyezm+pYhUbwYDqsYealnSoPJqrctjv5as9q9Eh9kBiPLxZF
+ra+5b6ma4oraofRfqvCGU2eF06MJbdm37oUduWcSfeCRXTBGC6ZnPujm8unmdRu
Hy0SwFW2te+YyQnxMxaZXaGt98taG6FLffTNlPXhYgAkMQeZ50HmuzEULzoeDPad
w3hGN9//ivFoJdmmJrydXCNwiMLgznBjNU9a8y7kikt9vQFOtM9fpJu8I8wupnri
G79PTGtZEsIZOwH/UOrWl3ZTNuUbVB+ZS/N7WEePv6hUAsg7DBhgiYaR6+qx1dn6
XUji8oUcnmH51VTbn/2z9zkhiXNjfh2cb8al8a9KIwwpz3o/Wx3XkeuDyH2KWaz3
PqFwAuVrS0MJJ5hxVKtJQJRWwo5ZacNNGTISow+h+JvDZxBV0PncKGsleD3J1RzM
DFDoo7e5LcDplGpD94V90VwGyIfA8Oj8Y5Zn3zjCZ4tugQ4tpJFfDG2K5pWSXXTU
5gaJZ1gspNaGgUFKYjGD6DuudgRwuqi0OhSVBAq12Dj6NG5ebKDtnwJiTlNzOHnn
RJtOy3wMOpsGIkJEtgy/1eFIXVR+LViEWQscfTOufGaEczKvF4pUCo2cPqn7W4pE
EaXZG+Qxu9Evutx8CzFhs5RBOaydy0tpmenqt/l0jo/F99MIWQtK31p8T0JU+pDZ
n/+UDi9OLWCx0ijlJ7kqrUUfmZ3+BUFkVZe1UWJODH1l4mZi1eHpDlPtUzeRKY/R
swPBkQRE9H+XR1kJ4ccfaSi/qFzzFy+BJko9uI9Dxq74nTdEgNULpcY4QkvoBShd
ObkmyWDI5SYevZ2TmRiSbluiiOGOZUNTYlScG9XYzGcN7YGvsRNixkIoS9A1vCJH
ZZiWdkp0/Kws13hUHJuOI+pw4qdd6Y8kEUZcncY7ZSX1B96jmdzOOkVBTjss4En/
tSjDvLfWeAyweL2wFiw3JGeOdz/FygcyToIJFNEWBfTGv7dDIHLLr9xfKyupjItk
e5c8jy7SEt1+yDQOKdmNDFuRIUAncZe0Ycw6KouLov2YdW/bhUTg+9SLRPh+2aFD
t7EH7F3Af28/pvpxRkF6DDhubAV9cbNSlTbCXO3Jg02VL133IGZ+Gxk/l+hiYbXz
lJSe+gYo2TSmg9Gy7WjlaxIy+3HGoXCr5Bpn/qbGV2C9cG9f2g66xziMAElJGzmD
hnDdtFF/HjyExYJIm1dNlu3juEYScy2Jfgs8/39doLcroCA8XxZViN1MdQJbsFWP
4A7CNz+hekPSy7TyCTTUIxcPGgkX8zhJtSjHZlvlURlybK630LkG93dm3WPLnAhf
jw0cHzbWMaFG3yyAGn+CMVEfH/fZxit4grnSKVXZXL7yzB4tvVbkWYBO9vKPfiWA
kd8lhlzS40bvnvOR+wLziOx+JuIutqNI03q2efrVHZlwvu6a5FWXaHPrkk8sM/FV
M3fQWtdQ+sT6d9MzDQWI4iqut4gXfUIAXheLcpyz6J02CAwMes74pYFaWBoyqN79
RHa194aRVMv19pfavb28abIEzruQWbN3N5EMLmvvwAYcWB2Pqbp/7J+7iWLroaFr
LBoqzi0f/P9vPdz+eNI3gWtTxeKLYdkU3eL0/t9jyYEklkGovP26qe1ZvN1KsZnh
UbIKKCPzqjaXBccEy1HBBS5Qc5Lwd+hlYIyV8JEzgI/tFi5MtOKMRup+HQymQIM0
x0OQotD/g2ZLujrVs12i6pZOuvewgs6f4vw+bLomAZYFtiU7MJGJVTT4rGAamILe
wyPN1+0aXyeX+L9i/G42GmwVpA+aYYiUkhWtwaGb97O5XT1HgWyzcxk1ERxKV9k2
uj0BUjPtJPTrKVpxW6nrpHs+7ybUGh7LHWq0FhZ5F7FA5jFeG0qmz/oYLNAq1T7s
WLjoEsDkfpaiqk88QwnBVgxBausdgIdo9D4sFVN8ZZBRLa07goTlPSGUahMtYKdt
Xw903P6jlp5ahJjEsTutEC3y0QDgcnC+bjuqq0yNQG5ou4ta29RurGLj8/Or3h1K
cqD+T3knwXTDbg2Wc3F3rlownHEpKaQrPtLR52+a/Ke8k9EkNpKWZ5n6XZPQJIwx
fWXs5L7MjZgNXg7uUJ3tEyxi9rGQbldLNLb1O7J7VnItyO5RQCwhxs5vhac5Soca
95ZD5aQZnfGD06zpMOHGX/+jHkWJdzMrmaUxvBOLwWFc/vMvcBfUW0egsuJwh8Bd
cnLEHFLnbdTm9c4BTamODtArT8DlGdfiElkVwaNa37fTpDY+Xm1hgYtHIpDl3gNE
FzWHj84kY5ds0jLv0O5iR4EI8w8/8GLz0RnQUAXFnAaKmATaX1DouVOFTe1M44BL
pkcM0+tyKBxM7gJaixb2twFNswfrhO8w3vm00kksbUT9bWiT+gleQ7+qU9CzJsmY
rFM3tXsUnV0d1h+IA8gcwJAkBsibZaEzYu7UKnwcjRqxb3TYFU7tsnIafVNzvmjV
sxvBMB1h9tO8jz4a4DiniUBWhHO6XNXgGBfsowJKUJ0Hl1W6fkU8/p3DCOmq5n6h
PFVHq5IJDcFf9PU5Bmnu6V9MYZKyM0Xz+UnlxDXDpdllDDu1KXkJa4qv0rihPt7y
spKgoLbCqwxtGhgH0qTgl5C8Q5vswmQpXlS+bisb4TAuYSekROza285+qU+CMGUS
rb9npYwB702H01hOnjUOxfxUD0VuBODvUzwTusEphFvWQGSb028v1g1CLQdDecwa
VTR7tp5hi61pKCfmN2dON61z/5ZFeM4jNeHohqvEUpV4gmwWr1cvhKWh1AFfJImK
LNPTWYX+iTXQq4ftZOh95zpc7q8ru1F/w22QuPnxTcoky99bdC5kxiSxpLWZLLA+
g4bzdD3FzVrXs0YczFsyp+pDX/mrv38R3YXcIBrblQYsDWmzXYIMUQqQ/nBVO6y9
sWBlkI9Uw2A/hJA9jGXYwch2D4XSHwV8VA5v6CzIsQFBTynYgzLpbKS1SsG/tqdZ
YiGI01k9tcf/aO7BjqiWkxjv8QTKkGOtkpd+o2IfO7ySI0TnbVIwP7VcFYIx0gV6
UNgCfu+6VNJt88wyHfYJkpxSAi6Bg35OvKrlSUvwAXqGpZYSW8/VmRZiZShc8GfA
/U17UWoVXZ53yff4X/ol3xK/LU5uNYbbo6EAy9QTcaut6uE1ArsC83+6ohcemTG8
28hVKrG60DuH6HQWuOliTz9Lu4F8EGFWin92SACQ9VCDWbS2dZYZaGbGFLqQy+cY
fm+0sWzPP+ZNzE3X4p2kRVhH9BmoqD2fe9Dzwc6K44g0Y44IK/apFHO/RuAreduY
ZtusCSuPLTjogp/Aw1NkQP+fMeQXQ+Yp+8PRUVBXenEqGdMakB06NCK6DG4f+SDB
n9KMJjoGbsw1pIl7O6MnsTk0EaKj/gs6zGPZ5Ta4pRUqDMoJuXKKPjc2j/mIJ9v5
DB8j9A/U1CZ33KMy9O7Des+qSegGBLwUPH4ZqUMm+gD/lqPacra5d6jxVRfwK7mL
8lw9YFIUs94HGSOZyZKUAV4I36Ns/sMu39sFUvg5t1oBNLhzJ52hvhj5/0pO9dis
cBNJQ5i0OF6BUCZuxK9xynbpiG6ghabWUaJq0X+SvxPfRUN3TYHyIdbqkG7OEV4h
9FMKxK9vFr3PSlpXeyvRL1Ora3E5yvRsQQYy3tGiaQkiLQgaukqNgRagf1+3GV27
W2Ny2Nllhz6NHiQSjYb/B/z8BBmAf8f2btTzCJn8W1NUX5DNYMY8GMowchwP7owJ
ZeWJkMNxtw1c0Qc2eQNxPwLWKb+MeACrUTJKgbiqiEkOFxRgpEvVtpoE84OcAFqa
zaMf4d5ZG5pE3iXQgRcLZjhM+EjecVwDkOBiYVtMwZgeWP9JA1pUtaTGTMJjE+nM
6w6xFkPdINydnuGdxAsMC6y2zjXokMKi0bkIEAUWkNMCPEU0pirCc5NP2sxhKf5t
K4AUPPKZ0Eigy9rUpVcLx6Hywgsq3/PpADZP5+rDxkecSIZd4BbtVRjHNMd/hqA0
p62itjUFfgblqSAlqi7B5DXgqhyKlt2s8BQv3HITtXl9uHTIUpP/r/dFUVhWMa6P
MkWYjWeKUMyUogQm5ihVT5eoIxnUgd55akMmBXOuycQZLjCoTeLFZs+G6aqS9NtU
9HF64dd5ThRXtO+QIEjw4UtJkycP7pGB1LgJ+FHnhriJD0L62LvgoPBJyOejyuf6
dfJA34HFL3ID98gxrpTjH67bKuNbFlkI3POZPqyIFILio5A4qliVHDfT2cxdB86R
M55Cfi8jYL1yP0XLuWNy6fGt0JOdjw01xR4irKJhKRXmhfhTv/luEfvTCexDbrkT
EvnWOHZpZENKLEOSJPIsU51HQQdo4x5QT+XzWj/xU28/QAeiTQWyUqgUqnk5SK9i
NmHJmdybcv9bx6tEAYm5DC7EWmQgE8DEitZag24EPpYzepZQxo0FM5hcliGz7g+o
3t2tL3pquHLAPo4QbzF3EOhqHarZo4fPX9hdvCsQMdbILafQ5osBlbZgmrboy9+E
81wOAzO2D2U+GduqyjIBfEG/wNA2ERPeNOMUi197IZuSgtAWwQbkNufpG3REqeqF
p99ccV5ZfHKLDBX4HYjQk+mdpCAGnf4hEQ0IEFGhRiwbCpDLqPjLO7esd9AUQ9ZF
Tdcd/eGG9G32HmI+bLQY1iUnqRpW7OlXjtZ8/s1pM2VcwciaymTxuyR6UoYseeN7
DTFxDp/tcFhFyKnyLtV8WBHG0SDSjTC4ncsZ66vZDhdr4VyMbUy5nDdipk9V0nqF
W6DBv9yg8cq8R4lBVe2zBRZjLf/MeFSXQRQS6KwgVqoS0swYlCa9IVF70Rt9YG+l
D82I37EePKlWz2ZrcHP6Fox5PmE81DgLQi3XjgEk1R0lNU2kLUBw+KI1RqjUacZJ
iWT5v3HmziSMPBKio4eqN+tX8A0wp6WnE5//BHRK75LUDXaU2mDV/aifCJLGQI8D
oRyNxgRcwv5sQpkur/A31GqNEF1dPtR7h5wed8PRHa+kc6FzltKn74mHrUX0pgVI
MmnMYQTJ8hwtLsDZODecZt+9MeRACF7kHbXVuZObbSfry6zWLc54q5uhXWWwy5Bu
Trcp7Re+1iFTL1drL1LnDDvdGJhFJwwh30i1IRxUkKZvTDfpsNmXOaglvRjaJ3vK
4K7BmiJPbOoR3ERf/HmLlP70DVl9sbSXowEkO5iQDvc4+uGiUYPICjij+PEHkY2d
sGWTFylNHdW1Rc6ZwYdCtv5jTyRzlAD9kW0TYuyBEpa+Kv5vGWnhWi8BXSSppPBp
e6/OTIGN8V5+VQCROqokk/T79LaWoP42wzZizzyuQpHZEN9vFljU44gEz19Cqzaq
40UuyX/YIPwXhQRydm6ICjlnMCVDucNylNHh3ykNq1YkBVpNyNW/1fhsGj68/stu
Pvc5xOcOZY1VotUgNAeUsZHicAoxbx9JgIe1XulLMM4T/SOtawZvAAvLTD4pvkOd
+AudxA8RoXQ0pHzp7jITV/y9Uf3A1wDhyMksmJ3jhnKr88YuOptICrCkEqg9e8XV
c3rL7dFdoP9oKaK3rrQoJ4n9PAGonCc8bLh4Wiy5M4bNZG1b2fETeQiEwcdQdSlV
GZSDNWzz2r6NUu+eJFXJmpGKumdNusTMfPU0l7p8T/Ra8Sun2fk6EpoYWaUEboBp
tsB7xRxrvvcLMryXjYrz876Wj17DE7cloxczfGa7xbU+agCV2ygxpocd9VI1sGrM
Z6R7KRUWqBP30jbIBeX3WAR8PbIZB3jCn100iefmnng7lhPg1a8VQahAIVgXhCvF
bAnzV7FSnCyRvRvOBMMt7+1bbovT0dW4OP1KUWr1gwprRxE5e+AgTBF65MO/jY+d
kiNjiiHPAK2b6P0T9oQtc9c9rWLK7r63plP31ZyZSMviS9Ge/jZ9t3x+HE5aXkns
cOICgqdFxI6yb6eqQF3qrg7+8+/uSwb/zMVzakih5NqJfJpIjHq3defV8E7YZMIx
1fqWUAu6XylqdJv8/25GGTmwAVvCpVSjDkvlhhoJvoF863NgoaWgvaMrz5nW+9gJ
n7Z/ypCEdLiAulFRPYmVq23wTP0FqME2x1MESlFoiaL4RCgBnfIcwrwjHDvNnqbf
T6XGJ0MDAFxwwo1ZeMz1YE1BFYv6b7jNoElpCunfRISLL/9U2PTqLdx4y1846SWo
ou6WW25xW8UNyGoalmVmDPxbSx52LuaONmA/In80UJUFEhMWTFJLgYSylyh6rfLY
G4YK6XzBbB3IeinzKAfKZyhUeR4G8x13lTlUN4Ty/p7OL5cOZ10Ea+uN42bfqhgY
Pnp1RbPaqsrQtl5A6WEkaMrtVDTJ+5o+6G+F28iq/fUcNX19qMORxmsGXCHLEUOB
zyyjd+x4ObW1o2BfIimM2TCA5ho8B423aAcyT3s+1MV9i4a88eHKZQsRU05ZGz41
kQtdpcqH0mtCs6UHevkU0GS6CCos3JJAtVUuGUTuaJBQfWfm6s7qifdx6A96P7XL
gSt9tLiwJoHoCjFNxJKscn9PxDQ0U7YAsThAY1Gnm6sjDMgCY3wFKBg9RWRIQtqi
5rTvCi9CedqMm9Cn2YyZ//tXJufnp0+U2+VdHNZVGZ8L5fgWXnWFu0Qej9hWz43R
/nyaVoVyWJjTSfJzZR5Q0kCq5POJrlspH0R1NZmd7dlPR0wAU1BWFWyqkLtIfxLI
qI8PgUJs8n40mZayHzbEiqykXFDaBopoi6uJkYBHhDaHNbjjdfsaG8vgTjSSbty5
YzO6LCx0SofhsRh9HVx/G+dFZDfYTHarPn0USjJbEnPcZOHOBsmJsvFaWZLaiigk
25R0AAxW3uMq3Bu2iI1L4Hy+NULv5ftAfznFoZa7EIfVJbrjHScKPqKdpqvPn4jz
gavYheN+9pMkgIbCRXstBXNFpQNCS/QCWbXnCKwWmqbTC/U9A8JF2FDHWhLbd0X/
of6vwzwZpskuoCtM0KTV6JxPJ0F8+m+BuhgF6FlzT1ajYUTDeoA+TRYBox8ubBtu
kdVwipS1tmUwadDwPjcuMJePsuSeZsEpHAemEcsx+0YXKJK7DJdTSzsY7Rwj6wf7
6k/ZKB9MIf1BPd1EHZ5VimkVQioUFByKceUL+7Y4YkvPkFJtMeMg0kLg5wyKuJKK
a7wQvyrbHxgAWB1gYIgSiedTL7MJcxTb1yRYE3rxFCYfVuy5rTzoUAgCB0/st32r
jLpxaM5PpjdPbrJeiqCFLqOJGUnSu3kK4BDhtypkFqnU5akJFOtEZ8Lo4uTCnXRZ
lpOsLCPXPzawzTzJTsPB7BXXkaEGeajsmuIto4aakimwywj/33tOJkIAYMG8D4RN
vlJEjUy2n/aiEF1HxkAvjCC2QrC/LxcD5zY1vLON9tMFPPc62Lb5POhgGp+vwVh3
hn8zV0qVSwlqGcDuJ6NTYihJuXzcAtbnqSpDOVE+DQwdQwnOaXj69/QDnVH9g0qg
wZbB/agdja7N1aFa+LvpFXD2wGogZ0iylw+GSH+S9QAtUewb4itUKcZRqjAoGQqQ
s16gAkfwYmOghnSp1+MMmpfvdxP/HOayFQSz01nYtNHgUhCSEnqmAOI5fLkpRfu+
Fuxvf5P6qYkREQOLaj22ha7DWF59L6+oCNgR0WCkOqsC0zDVXTstHE2WhClWGFaf
nmQszckzDqJJZQZmgSWXHSdNVKCOuVfn2TTdmiOOcEkgb3yC1Uowe3gFqMnfEowV
4P7Uw8mRMuWvibiBdvTHoIqNcNW8Ja94kQ8SJxFDB6+hw8wTb05X/ZfwSJ+Z9ggQ
odJ3AqeA4sWBKyp9v2kiWarAmMBk7KOFIAQgRGO2ZkO8kcsB8J84OhRqNLzBjiiq
S40wAt1Yj2OKrKQKNhr/LWkA5NVqyCM9voRuyZDAORrc22IA2FBQ7az4pK3HYT3o
cNdNkfGvwbYeY3ZgNupwc3F8gqoHt1bJcSpbFQZbRilCgYZvAm6I+v4xkfJ9G7Gp
2C8992uW2gSfqAs0uHsZymOyZdckAlbXHDniC9Ue+E5HvYZTeXnVulLW82ZCK/TU
CPpSQIVHzluqyj4NPYKdsrCS1kN14/mYhJsHjjqtcamEKc2fnpMnYUjo/F4LAwj3
PI/BW8kwjLn/s1MgDgmgK/mYBB0rGZjZxMdCthoFL7MjR/4IkzSddeDCPOI0Tbyl
RwxoOewZOzJsGTbAd9jMXnjQGxF4CaPDiLhHQjnRnhSUDerpNaV0iZJHYlgOSL7e
a3Pf+qa5yFTLUpuP41psPYBm4gdd8j3sgiJGqejZTze0o19z4VeFlPFsgMDg/dpX
421VM74oCGCW2ocpqwwnz2D/p67Ek3cQ+wyRlVuU4gu8g7OktlhwuNViosHV3WRW
z+Iq+STW1aK6Ir7gQ1tYR0Azs6Y9EGHiYddn1qmVPgqSjXECmUGynHXVMxDn6Wx9
nCTGnE7L2CesmNOqwbdlIoEm+zAQ4oy2lj8mr1QIADbNs62kTQKg7mbjEbAvqz8K
2hURyN27/OHf+7VCso3bSCE+/G4+jx/m18h8eKa5mnhBhl1RNBNsbo9Qzw9acpHW
AnUWEXzFhyGR4I6Z/YaxD0t0jWiQyBcENksA+Db03HyZRas4wq+GMx5ibdgL5KDR
1+5IIuVGJvPDCA9VM/LwTUKEDsZ9+8N4QDUAVixgQs/eYi/pc+sL49ikMJ3XuRFH
k9OmvNHOPrC7Q42YC3AWsJEi+5HjTjU1/G8gpcUnIdLjN8Ut+wd8DkyN5X6qVZv2
252HtTG4qfppWF2LeHUs+cGqWvnIHpStoejgaxCJrYa+CjxOhGHwjQle1B63ufPe
h6fXniYLsjUO48FIaaIje5E/WR6uGmOlNNMEvS8BiP0yaiLqP3x09AMKRtOYwHTQ
a5/X+PAvtzyqIuE+ZjWgQyyXoVXebH9C9e4yPOuU85bkw41QzRIB68TqRL6n2kKU
vNKW/VitLXt/u9fk+ySrjYlWmYjmVrsrUrUFvbq+p5YOjkzpby3InR6yJ613Dune
eFP7SPNVr4Di2kINiCNBT5qHMHFQ/DL3Wvk7Rh48NAk8yyus8yr+PhV/tkMaPkei
yPpNkaccfgYIMZ7A+Llw6owgSh/y6OU6D3TzXHekyHRrauilHf4Eqkl3EcS92N93
I0dcWEGZRqColBIETUUNDCUceZbhVJbnHZL5vMmmPno2n+kd4zMQ9d6EwzZCx8yg
dvFlK0LcGR39xh0FGeb48LkKYeAid2FB6UgYFsaFcfxuT0EaTFhe6TBOYf+PlgFI
PU/Qyvb4lvqsW6o20lOAV4rWLL/RWArCgOydDxn0Yi1aJQI9T1lo96buit9Uc2f7
sutLat+dOwTdzDvb7a52CSGViXE7beKSnctqxfp2eiUEPIcQzjOR5/EqsOytVvPR
ku+VNMO3gOFuP+Q7t+pfdbKH0lVek+d15Oh2n8t3zznZeR0Vrlu8mvpYMrdu9HDy
zdQBoduAlbN9xFC9mMs+xP+efvp1Qzpx+kdU1LSRBshnTzG8bop/CqfgbUatLVzL
/gpbzLt0DlWDUyIXmkngSCe9QADuEDgciWgGxMMDjHkmwa5jHlhqDWGlH3iJHEG2
vdQQikDUmv0eK6oO1tmKDBErDfHP/RG16OKO4Jf5j3xavHxa4WCsd7PtztnjCBT6
KQzlVBu6XSD1/MNFSoY1DUmfPOp4z6emwwnT1tKLZqkXoxJDw3wMKj+CdLnST+Ti
2B3aH5JVdFwS0iEmIGs+g4V6gf5/eMRKacMKaOTZQ2bgeMJYBlhQAFiTHk5Yo2DI
Lg7mDUl6qq33Dfvs3Z5gT5G1yLQOfXvjFncn8vZmgwl2Mg8wJtxdSSOF0cu6/xyj
Z2Ixtj6cPk4tbkoYciXm5duUgnLYyMo9stTj/Itk3MpEUAejtzM4jRPaB5oZlIVa
FYatqym5uwkSZ0Wpr4f6TXQcRjH3f7/3chBfVSJRSZ7m+bvTz5ZHzC+0W7p9zMWj
o2JKNPVriarfFQOGSpjXPP7G9clH+S7o4VnUZcmHSf2KECm6i9QNOz5su63k1/pC
UYbVzFUo+9IT5K0EVk4qjG4R7y2nt1DzgPXF0vhJGy8sLdLJJFS8SJHNsRoZM8H6
PfK9m1MPP5CRHaT9RVql+5C7Z/lSQYcEAWWKefxrUoRdvQvOABfbgYx4Y1Lh8oPu
Q+QiinZ27jY8qU3qgcGLDw0WtX+9ixy90nA07PkiCj3na+jcAX7N2aGQ2OzJWOHk
C6+bMquFCSoNGTZ2LfbBcJ8zmL2DX69jERButF61GHiXX0v+9JItgCPuHU8mLimn
YHyam6I0h7VIZgvQkj/cCD8N2NkaPXiUHgANGUT2USfPUWMVHGB1ULenOqegcmQ7
p12UZPtWJfQ9WPnyl7uDsWq8ETYVMNVAGd7ZB2WUYckqeZ++EU1RraEyMCB2m7Zp
/NG9qGSbhRl+l3rHW4BWX/r1Hf0S5kaeKnX5mIr5yUGgmBI1y0d2jK8hNWHh1m9i
JJjwvAb7mgjLo3ik+fCJ89iCf1apC0cDxEaxeMR5EYUL9NvuWXbnALxuqXvM3swJ
J+BbhsecFh1gEQriAPEhG9ZDkh4/Q+0C6Ezv3D8kSeMXy5S7bQDh/VKWcQqMFxrF
AqO29/QM1ANPTWNKvM0vhwv4m6GsskJtKJ68fE5ydECBp2Er7ZhJIkqgR1GRo1Nv
2A8MncllkbFy7dvb6wVTBK9cGBVA5Cq8G33ZTNgf++X21kkgY5VLI0K8lyJqKC95
sWkWuW4tZISqMRjXdlOucwu3S6OzVM/cP2hTQUArFnY6QoBceHphY1BHi2SjPD04
Ax9Nw2/pLDBlkS1+QWdHzyGOZ9ZzrdUk1SdZEBMI02HeCrNhpWuW2VNtn2hlq3gL
irZlZOb2UbNe7SVx8X6MHSWD+oMHAEgrvZxr0SOeu6hJlS8ntOMQGCKJDw8CmZ+d
XoV1gkYiRBqISqTXC46pvFeI+7awJsuOXvDBWnBETAA3ss02rEVeoNoqM5lie6Ep
Y9fZgTnlevWqL8tsA0GLZ+BdWAHsdBS0SRIQ70LWNPC0x5gmNEXbqDhDVdAFv2T0
kcjx/SrmIcznso4JvU4AurF6QfwyvOBE9oD2aFKoYVlx/dkhZrgh0YvjrtEYRwN7
eQpIFbgjyp3uH6T4EyFI64dm4+Ex+nFsHeHO453OX6EDC6is/2jCeCjhSFsMQgNI
dpBoxlCrn7FfAOqvqURX0HIPMeDBRAyvYiYJ1YaicxkU+uO4DsZeCpXSM45rdZSD
H7FqZzmsVmJr3IkddSEdG9X7PyunkWcoaBpbBXIQZ6/VNDKlLqj9DsgTUwZJpayg
LQ87pytI7BJOqv280anNkWe3i/DXypgnUU8Lq4Sw1tphUQwzhPuAp/Y4bNnnpgL0
9C99SRrwXpZAnRU/g1rIfUVmx4STEx4RBCc8QGRqXXR++agovRSfV5aR5qdrB/JL
GKlhmSvHa/PWCk1psWTNOp2sgZlxRFgn7+m5vBiwIVwFzlesbV6QV/AV4r0Sjc5P
qzoNcNdV71lqh3uUFphJ4IYCRBtmGdHFy7OJ1O+E7v0Hswp6rV5ZDjstOATNk+AG
7/qOvy7aZ0wHlA//35PvIbXj48FpJEtpp6yohxf2Crb5udW+bxy21XfpXsd1+ao4
1CvcKqVZTieqW6DxmeqJW7QFTsTJGuY1cAlg5sPTJqpcksLpYedH0MiA9gjnkxnQ
mGENKEzXMGcQReUdgpEjBKEIyCDt2hbHejf2rS7hlHdQORhoMI6pqCthEL5wwldG
hR0KEttpVS6ixR6n0AnwTcqdHwuUUyELXRxcvY9n3O8NVifDAHZVGD2o8nsyyO0+
GeXLZtuTVS/vPCVCSmo2rjiyQ0gbzYn0OrQdKS1rvHPgl624d2DPVFuL85X95r8q
Fo7G15UKjCcARGF9dJ/pyj8bGvVGTA8KNxQFWKRNrNGSvCmL5SHc/67ekj88+zGf
xV6jbyDUw98UU9eV2AmqFt2Heo8MUpk6BaKAjus+orJSzA0TiIEA3n4azRK6HzI2
rIkdo/Y6V1drvmKlawQHBFFHLpIVtRJEHv49NgQTNbIDfwIYELcB+fYcf4QVTb2M
HDGRC7+g642yA0Vx9Z3uM+CRk12wYu6LiaZf9W+V01k7/dapY7mZIknmhZrPd2hA
8BEZI1LJuSYel/qX1RvEhc8EQkQD9qAizRuc7qDAqAihSzZHiVj2hfCIpQ6HMj5R
cpBsqDH0igwv5EfAwYv36DBuenmbJGlOxwXR5YnGe3+jyJWoSJctg/kaYYukaKCy
wjxXOZ/Ys9uCTD1ZWXwaf0UeUG+dki0Eyshsl+hmxYHYNAWSDMBcEF5bxyEcNkHG
oYiKB6NKHwLTJdO8V+FTyCMNlA4juxX5x/Ch6PNQcEkSLxLCV/vLOXaihwx7Egre
ZDb48ghbkcJmovdeiEazQ4DpmtOAqT4qWCibrOMY7MaBVYOe99b4wc171FNj4ePk
bTiMI7JwSZ7yfmTqM7UQX6y2YPetVLc3ibrcBUFrdgPGWSdVI0eLBfL/JgSzV30L
PWo82QS3RnACTvqMg2bRMdapoShyZprj6TiosDocqUvxrTjGrLAaLG5G0XSZpo2U
HMOwKoRgQpjNRZWT4MCFRLLpxPx67iq9WctTY0P3IReZ3yDTUETHQ6TL9b4M18Vg
IwqitzrIVW1xoIE+Ymh3Kd6OyVqZjKTLgL48nHKgmbXJa0BCVAfKAlrLzlh4JoDB
DTu1GRJ5wvCh9TgCNNoAEowlKgeYcrOeDnuUUrTlARRzVmq05t5BY6jJDwCAqHfw
yq/7lW4UQe8VTfqpH8ocW+xaRezivVPY46+LksiPGCUqGPjQ4v5DdQGAED2b+ToQ
mRBxI6V91YmKAHQABs78ZRmlxWgsZVFmSSAlekK7Cds4Y2A13L1texlnodIkajNF
vQIJEQBGMr5RMYGTKq6bGF0HToZ+VY7ASTW+v1c0ib5BMzqVsrcjKeu6xbwPP7ox
P4TrOGyoh7kMpdQZr9Sh6NJYYXGp5lNWlk50vnFtDHl9K8b+ZJXwdTdDHSFeZsqw
Acie/pjrDZgZU1SCUxDTqCHm+/erlNKaxoToO2UQmA5VU4fMtrNc0GEpa7o27r6n
67EB+1rU7tckO1k8XHgx6r5dAJPeTCyd/SxVFZ+RAf9CRMwqykARZKXfSDM9MNiT
2DURbmiby3sKbtxR6nRVwxh80qrzgmbP4THl9c0mJMICiQLEk/QdWk+uiHOdWI0c
sVqB9RkEA63WttCyH3yz8DrVZxSTh+toCApMw2DEy3PdNrmUOLqMz8qnOMjiaSBc
FpmOmgAWXpxYRjz0alZar79BPaaTX9O49sIRlO+YGTfmkeFux8JYuIgZ4pRXPZjx
TYauJSx3zZAmcpMgdCxUbOyCh4xBIkQIU5c4cxyW11NX+rfZd3vLsflzGBvXhJRK
OVZ88RdA8b61ChMB0XAzrIa5P9NKiNKszGk0hFR7VdQFcE+Q7W3H7r9K33q7iqmw
RPLLBLn+URJbVmpV2BqjRIOJrRNAsqnZDSHgfBGcfOLtzOLk7wZj1KKLtlQaauj3
hTWUVSDAldDiLKYEG/WmJs2kPNxkuCfbop7t4lMVpHeOsOQtxXRYer8W8iHQaKw4
YdYdPpZUY28USD8NsBLtqyk9D6nebQr4KDNjbhlRWpK35pjsLagX9FZd2P8d7wlU
Us64fMvXx/1QDzT8MlAs/I8MOms0kWtWJfzd71DBd7+7EQ7YtQgOxB+pigHbOX/o
BTID4nGX+PUyzm/cuObi21bM7aoJgT1oHdmH+dvc6V/o9HD0jiCXI+vxUe5fdzN4
fd5O5LtpCyNeuQMDFvgsKr/HDt1N3COnFevJJDDogb29oWnD+Dnueb1BaUM1ICOf
hMQwt+ppSKmzsKd5YATwryv9APr/+giXcvHMq+fJhyTQdtKOrDaw7PK0IJnafwO3
V3hlScKfyWn2ZTAhIBMqJ6xE0wEFfOUoVLh6j3lmvpKEvTZ3TIWLjBtS1f4QJswv
WaDvFhFxPBzAmkYofYULK86nv0XYtHkt0HJQLoHGq5l6NPc1LTyBxXn2bUp1tPn9
B2xrdc35mVELcAVLFncpOTlnCwjYir19N6TqS5JPqvlDlQMfnBOhwHRjehSCIdPX
UN3trkOk87SmIZU3AQ+0TEYezrJM491nj1w/ucedwEoY9OFJ7GjbpUdecrg1kocj
W1kAIcYSA3w9o0s8vkcDT3j97KL7JPOBsnTcch35rexuvrztq6bxBo79C0392OW3
gImhhc43O+QjqkyDD2NJJKOyVB91XmCCtH70FL9tr/CcfCpZJj4jBux7sK1U0E5i
KSKy7qayNzxDr4QLlmHC2qMBheQQHhPZ8iu6yagmoFyVFCfNZE/L/O7FUMCUdGHC
xwPNoxaFwiDqyZMTblwb2fMUK7/trz4nOWsrhbE4VCw06mmqiDzCF/y90dLcMIuS
AZ87/9BDstDjfsCQS5oz3g7yrrAjiOPLZ21hN1EFV2LurH+PeB1qrEPJjNADkt5q
SysC1/vvhNCWQ1Jpk0M8omW0vpdM9Uu2HZDyAQUbX1+jtr/Sf5b1t53RsT/taK3y
faKDWqjEairR+Z+jxB9zWFmzmBZUlQCrehRn0lAARfm81VUonehOMxHxMyoWUcYk
rWFHe6pgdZ74AI/MD3oeB7qxXvnSfBombzez74m9ekO9vl7kasoD3giEJ8H/qzaG
KP+05KKSidGAamyO6h/GYFmToUjdiZuY0iat6iZYKfVqSe/7DTLhZ1W81ySAPnqW
a1We5TvowWOCwVEM8y0M8XOCZBkeg+OlqNIEeev/eQjIrJSXVTS5NNgOJiFsZAWD
/FxFawpq/rXqQqa/hImhS7R7btkkhbxaPrDiY4F5ENZmH00griByA8POTBiHkQEU
gV40xWrsDPgdbrO9+ZzJXH0ttv/RTp/V1EPIaOR8/pgtGbI2IR4O5OHbzsije1zo
3F3/L5RBBw7gUn2JRrKbfRe2QLpekZkYHH+b8+GkyCLDUDetPlHrA7KWxkhx+Il0
G4N+bg6MxKUJXsY6QeEJBrGic25L7ANZfLJK4IwrncpTA7T8i2wNiyqDh6S6at38
mSURTY2SLw9PrWT3yNbdRWU1Qadn7Or32O26rz4pN8QyrEvng6aEkW6f4+K/FH7f
+WY7ECZ9RkLVUUtUw5AdwIHiyRiRPTMp8QR8dxPRaI1mgJFmqTYRV7CWMRu5t0Zy
BZGp9yzvuHcNtG6c8gN/Q1y/zjSY7WRjnRlcRgJdvhbGM7i8wM2KvTIGXBIc8JhP
WWqNSx/TKZwkYTZTSy3mM6MrS4m1lay/7gSqFPhfzGNY2UMRC+/3qmJ2awcIcvNS
neFnB3Ri2unv3Xef+kmAAfPZUQwLM+UaKSfxgMIBvP0pDT38nRwNKp7Mzwywrij6
7qTsUkKCsN6Yxr33rVOvoLVmvVNB+FpPKoz/SuRxpb0GkbHxUmVYkc6RbG2tsXC1
hwP/6XrPwP1+1CcM9BRxs856CBzH8ooccuhVnnp7F6fUImHi+8QrZKu4k08auGSu
JqwxfvBOqYU1II8bg6yfCGMFX5vlH8NwfdT1i6BXoU5tcTIgIkLUJlJM4h9Ew8pH
KfuHFTxNPXBGvqduZ9rmlSvktzVzavZAD3kKeZtNKdupbakLeP+J5uqtLmbjdIBg
NSJrSRbLkpSpxn1OOBERyVfHl44ROpsluwL3TxyHu56T1eaZr1gSDbWO0XL5tdbP
gM3hk2cozBjiiRk5Cmlvydrt7CgV4hL9t4dUFX8OX1s+ZmosqPlxAGccOta+jUZu
tn/vhPXxYgJuyO7W35bhPxRGeZ/7GwAy4LUQ3FI4VbcbKEOneiFzmMeu9kddMDRJ
CiqE8wvorSAh49gvUq0uo0k0BbsAnN/EvYPMIInrJ9FM9pH5DCm7qdL8ewMMPNW3
xIFyK2US30GRrrMCDT7HnVYr+Ovyv1fC8GQAB68zeWGbdThPb//UhZZfdMRhFHAh
/e8H4xL8d7JWRjZ+EPMJmMtS6kbS6XoeeI5/R2WiXtcK0/buyRfjugSkmCuUbupU
n1UpS61nKoerv8ZldZEw7QXCLenAN7Vw2V2f5kQIoiUD2o0vR3sscl9MREjdkD68
U2qkQ8cDPo7JAUJzX8Wn/lYh/VDDfaD0om+CDzC52/fJYQbGY1EVizLdtdDGdTOw
+m63s0HYMCmMVIPF4JNQBXJ6nIyYQITwaqAbKL42TiZn5mUa5mK/XyxDzi/puqDD
G+P5n034+6Bn7udTG0EcqRk5VjNHOQDxpsZmNdUJt3wOwSPEJ9GlYV4LX24Du3pM
s5LbwukMvmRuqUatg7tT5OdsSOgJeTi4Nz4l3STPf8UTv+qtE03s7mspGUtFqjlv
4H4/aVujwf0zUdSnCH4L1Z+uJ91UxI3S3CZ06/aO8J+U629qDwAi/qMSoK7nlGBh
+RWLZwegO1pTo1zw/FR7zMiFf5EMu93u4KruOTrUiB28hR/Xekf5rpM9SR1t8NQ2
JSStJe/z49m8DFXtCdFSZciDt98VhbFkW43aRxir3JuZ3abt7LP4Gwqjp025kZEe
GtzdzSrfGXFM6CZKogBfchlWG4PIMJkRiAat6yM7yRiYl2MarHagEu8GiH9FuNcO
O2MewYE8W6ijs3GQg6M73tLv8RAZiR001kNot5b4ZpCBbDCy0Gl0+6stHrZ+HeRx
iBtkPyQgvDP9Rzwk29aujZ1OSb+lqo2ciaUBvKahtUJOvjzQLvQ8p9zNBydGWwvn
EjgI46lSJZ+NCiAxC82nX8BFb1geZgLsH/FcAQi9A7kyMA6a3719E1o6rN54Ehog
Z8TOFi2bCyJq+8j81HkK7we07qMFaBsXUZSTd0zejz/4IQbQD5u8daBr1/J7l53Q
Qh4bN1qrpogtpmeT95OsCol0p9npVAx6zQlz50ugIkOX42aNdKnB5SeAiFZalFEe
ToyA+nctb6aljDZ19sM+4ocZuNzdbczWz8v+KCehqD0vzYjyKIaHcsypNrUc3kZH
0VknYu73urGnl9+VD2/AbKC9I/7rB34Bu/Lo3ns3yTrJqdXx3MKOK+YfzI5cNRbr
41SoaFXXw9mSZ9vhCl67LL8vsEUqfZMyNHySK8d+vPKg/YOEsKOxJ1BPxa69BUKb
cIbTwxqIhsiDGVxgYTHPQwL3Q/CHRkB9qPp6hpY4J6Ol1DocBzR/T2PS58HNFnHH
qog1uaxw44aPvUSvtGzew3LyXoHG7WblPnPvml+AvwwESg1ap9tPbyaPp6+9J0gZ
xrabqCePWrhQzKM/NP6uRnhzglK6pfSrfOigHihfU/7L/o8eDvnzvjJniYGupxpb
PkCiXgXXcVOuCFoUyk+Kz7KP+ILhTos4b/u12RxS7elAfDxD507zwqMzRdAwhU+1
eYvBtMtl/V8AXmIJpnxF4ZFfEI0eB22Va3DqBhQ0hPeU9Hsz4mXFOD47iII52nAN
0LiyVRjrL6GK27NiGwrmWLd0wPbZyblBlAsPkAElrDgOGdwuyhbn2bl3Y1s7I3JL
xLtxW1knKKfq4FTNNtwt27tF5Gwk0gIXukJO//jsr6aLGxb7wT/8kHkDG15VhUal
shye/rpHJRe3hrM3+9YUut/JeVlagnTSi4O7YISXzZty8LvZpoLlZIJ67pf78ABg
Ihs5OZWHhdIO545JPEgMy3Ij3WrVHXVlcxzDWvfD07df++WoymXaLSYTq4uMHaSL
gwCF2chpb74sDu2eYOx34D9kgsMAcPZkvtqdJTekxFUI3HMV0ghjrJykY3a8Yzwd
VLpX4zKfB1JZ2t7vjo/K+4WPN9qUg787Pn6rW/N2jm/2DPc9a2EDs+vIEcQlVG2C
b8mqHciNXl2D6Lsaz8L94o6qpr2SCXy5RTEhOm/vyWKgOEUDexylZQR4SNIdkRyP
8lQdq7OCT97uMRX4HVEMd5pbNAJopMcaU1ue1whZyPYZ8daNzvx74KszHtVibk9r
eHABzgtf5b8DjLgsNMvXwg5Q/eAgCfurYRUw56m1UnapiaSlL66/+eQiR3rdw8sQ
07Y9aoQ34fK2aozc2FbFpEDuAU5vd+WqUgvl6q1uha864K8hVlWlGZfEEg+bWCby
u65TCDmZwKkzYsA71u03DWp2AA1klSCamhqqrbs6xhVQ2Q3x7mCFomVz7CQuG+Vs
L5bh1OES6LzbD1f6C+KjZ6pmW8TU4MeFqepJ7iKWoBArmlnwqu/ALiWenzzj7pTz
x2NN61mUnsnFMRPNEFIjTsioPeLZA6hM4nnYiWzmgTJKo6bUp6xyPJlZ524hmwVb
+BnWIj+Wk9hWuU5E/2aCny5uVyEve4RaR9D07dYtJ1DFGsFaSNlATeOmeuapZa5n
kV75B0c8Lsj17C4CluIiTOvMmgkJNeznglTyR5rfBCq2zCn1qTeVx0AhsL6YoOvy
1jGF1KgWhrwBoxxEDStPZ4MeVBb5iRgtHxuAb701L1mlRyKx6//7xbp7OTCpXHO7
+wh8YmNY5l5ize+hE1jUQX4wBq72h3j5aCGmdPDUBsKzXrNk1KIPvIRG35Q7lQ/w
WtpFphsxv+OmWVm9kzfkNtlEuBC2MxoMnNVnWFUX5eJFlW0DRQbWY3ov4h5VdkV/
NCglh9GTZNBnngyAtKPg+3xpFau09agQfzth6AOMcSZ1HcSpVDqaYKTsT0/IwQR5
swUqDDfWF1o4WKWsurAmsIR4zkTl0/FVhPE/JuEB8ljSGKw38/qIYt1Z/rnO1S1g
plfSb1ZOOYlQsk5tyqXsEIimZARCbo2V7GWzqb5IbLRxkEypZm419mfQEOPp8pDh
c7BrdjF5NBfiDq6Dhbh11eAt4/OGAcNrkfn9ylH28GtsTSneqFQIWXpEFWMhYpYs
x/rS68IyragQPphLVmB8JcWGVvtuU35jSEafuhCGx6Wpx1J9X84dmFGoWF1OVWDP
ZDQ7C5KP8/VVi889FpHlNbd5x0ARO2RtEUQVFwK6QpsifhORv15JWTZeJJHPwp2C
Hr3amkFcBG73zM9EFw/zrihzFb9iVN8eADhU6v0zu2ZZ4Q6WyE7dEujzxoJyg6vY
hzZf/nSVfAfz4XucfbHMwSpNbgo/5tjmurFNY88LBNkpQRZNLeoBEMi4F4EsUIOt
T2o3UAINiSEGFju8q4B45ZkCSJ0+BpDtQM07SIIKHJpiFldt2lRboivDveO8GSzm
w5dNeFjy8fT8dAoC38zSyEqan2+VtXE/VNsOvVTPXPv5tcK6zPdi+78uWsNWaOtd
2EeyZfG5E/v2EU33WTVFxjZ7l+HknxddoI6FAKodgVGpHz1Ce6hNsGdEBFuwZuj2
eK35OqkADv4fkIsG8tzC+rIQnAPIftuxySu0/VEJzuFo/R1eb4qTCSjNxabc4I0H
p9bx6k1xdh1FUrCHNQN3irPNiaF2FJuEoiI1n7MFUE0Vvym89YvaNuonTZeJKkqK
A3Js65qvqzQgDmjQOBn1sC2J1sJiqrnsR+xAtp8+/5wA+/FRTyxiiAfPOvh1k3b7
mGZTgW4/ikNmWfi2rqddyBves5/1+KfMjXgsd8ie4xUZ7rnKCwbqvPdNQOwvQN2O
VXPTFMhYtuL+NGb6LoAWvGMVoxhMpws2K0nwQunLaN9+0iTBXkJmkuHlHFsZozei
9cNe8VGvSmpOuj+amUh1vDfEgPS9s7iAeg7myQS7iEepbEJnp1pxLMZGMgNSmYQY
Vxr3PxSRHj6VbwfEUjZCLSmzPdOk7t/EJpNCH2ly7APBZyUMVpqJAUDCd1m0IhPt
semTXyy1sybVivvm/F7DV+ucuAmmztMDFGnWG0uRRdnCG+IJh5Tf+DXZmdvcIEB0
nh9lt3lqhbKJdXJGt9LNI9RmiyBKLTIgDnt6FHFnx+CuUTZJkYNqym0lTTB0K0kW
BKT6rrm9FxJ+p5e9zsXSB5UoqBrHa0ZYQ6DabIPyZID6US2+WN7OGBTpENOQBLq2
9dqE+NAEOmsig7Yrs/GGNOjViu7NAIDWyMDW58S4lC2d/ckRGOj1oeoYUSrDfqP6
BEbB5jw5dVrLSHoAo+bRRx70MRVP94Q8o4rY2fV2QabpxzL//AGSNC/lLrRUkf+/
aRJGnHOHN45RiX0sE/mmERczT1xerIYWZPww5d6iWX6MMrAc/W2gy3Zsws4iDDCy
NZd2UVcQ1S6o7YXU12y1vE8FfF+kc2ZN5Csu3XODaYu6lx2bbER4v/GAzZNsDtGB
ghn5aWXcxrW0jSX6xz3gZmp9UlQiyRu3/ZLeY5p4dhWgVcrUoJLuuvulYbuN1+g1
Xld29QQCNBzzAW+g6H6ki53NeP6Kj6KWlpMonoXZntkKOti0Ds0Qrxv5EayOLAuS
jYGurc/ZrUX7+YdfZle1MMLk5jqAISxytZOAMOP5OMI4RFsIluiEUXReSIIr4jLl
IrCRSqeiMFrN7t4W1dv1tr+nvslpHatobg+dB2KNNuz2gXQ80RURS53S7wU2wde6
4h1/gu2gxp+N3bRkAYf8WUgk4CQHtw7DHErUyevNfiQwb3zXm93TQclEoBnXHu29
8rj4Q17Q8WzYeIOPB7BAAqKnoA5XVB3aJv8K2HVlzw2/FNp21qfTLlIUFAA7prOn
fumZhJdnK8vhGDiGVWUK91ikzr3JEB/JztUgyDy6eYhcWayGNsXUlFTvx/Ne1gYF
vRbfPeJ3Mcxqq9QK39KZpdbUqmn+H4M7g5jA6ScOEVj9fB6tnOLPp3nl/CbluCQX
lTq6QD7D68QZb6Q9bjkMGyx7bAUlvUigcS/3pIynjv2ArOe1mpoq76kB3tYGz8Kn
oYY5x2j4VEZMS4DVpDxO1DSTPgARaSYH8Hbf+AG9FdBLXw+zyktD0Y6m1n2CidJ9
2RFxaTI6IYcjoFLi+JH6/UpzqAH++WVfxw8OvgZUCNhORnwpLIXkP+eyOcEb8w4J
+il/WrFwlMb1YxZGXsxg8v4wKXqk6yL7fae72jgxfzGNFij2YVIMeLdQH3+34mAG
4ga3qxwbVzFfJs8GX+/C6ny8PLS6mMsTmcHxM4VvRdCEmjqUO4PyDufzDAxQ9pE0
IzngrbfwrdM1qrLh42G6FvbXvGXqKQ0rzyscq7PSqJALpsJ6tLjVV2uYeMlzjgV+
qrEhzJJ7FS9H9/pC1D3mtTwpyOLrG0C0WfS3aK43Bqth/mbnPy5q+dXJOBODfFvf
qulg0kOoXpxdpk/BlZEMTcD5J46sejmYyas5+7p2gsspoxbUU61fhf7r9EKWF3HZ
S4pHUTwUlC7JarDwSkxjtl15g7rY4qrJRDv0sWvPWlZUEFw6Mt++ywIYs7rIWGPQ
vUghwrIihv/xLDGww8Ak+yYJcx2Q8dz7aZaJKm7qd+bCTsOXR5PXMWQ4K4F6a4GF
YeUDGrlNqDCrcKabzOm+p9RQ+XJ5VQcavwFiH5Uy17F74vWwaGbQC8zrnfuqLQyU
02iLsI9A8CLQxOIrwuHHUANknkSARgcoFeMdHKTvnkLcBmy+RalPzKH2PMwp2dab
aTA5FJLcP5B4zQLThkKX+PS3NkSrn9FyBMFIYtJV3bpdjuuefgzUzWtQ+JiYCycp
DIJoZByYJqgwKqTumLVcYgdmAKbjCSoJmByY1B1x/8FpnueuBTXoNsJWOXtysZ4n
/8rKVYluwkS2SHSRzSlrRGLcf9Jquu+//JkJYrsN/JevAUHeTeTdo7rFvSY8pzUD
J6EysyJZzp3tbalU0h1EQU/k40mFMPWpaUhg0rKmDpXFhQTgkJ7GQncbfH0z/8yL
aN8/zzWHCbuDv/glDGhAhVVVqlwMIWnSIS8JEoLkh13jO0Ei+hJlbVPyH78iVMjM
qchNyEM8Pq+58y32R/4aNCTC4wLhhCyJuHEBu+fbFcBZH5JtEoD/IumYD24OiF2N
cemitPxvCUEbyY8ZqXbpL5nzdeh9b+G2HV6SB2S0dnOEsrKnfkoSK8O23KDhacE9
1MWMNmIOmkU6APH8PR/+a2v5R1xo5GDl8Jj6W53PJmZyFS9dlnFgyBwwLNIWBkyx
TohHtKx9H+Fag+zFrsuN2CFkkPAG/23Qgkyr/9VQvCUd2zum8CfnmTkED2zNh3vA
RkTNM96V+04VNSLMsX5S2Xzc4skNoehngMPRtPyRDBbyQAsjvtw1IK3oo1H1JQY3
7IXjqL/omUpjhKaCSGe155rrx/Osemu4AsGHL+d7YEDoYtpdg+HiKPaACBLMjcu3
34vAM5/CGl0p6jHpKMBqb2nLOF5vBB6LSKXQ/Dhl9eTAbsSfW6dObJQ9LZ8bCI1D
aqZVsHjMvZ3arrHZ1s2eyY63/FdY+er/xJ2h8G0EdDARZQ6+olC3pqxnHpZyCwaV
F6hk47Vh08XDrPbZmLJPCeA0ymYqLyiVvZ4l/kFaiUxAeCQTn+BORU4MRxcE0w/u
m+yHlvhoerupcgim4NJSDiIsijbxnMU3sy1LHUpBdjpcUAllolwEbLZ/1lt9c/cx
Ml/7/UDCIpdQmwo4P+EBAkYgAwjUEpwDAf9Wsi1kdJWAQl2N0FYWyw0uD7CAUOHx
VHxN3V269RTk8ZT0gJ6oZUBAyi9PDiVH+bNUj9Gwtc5BAITq46cTG4O2FYsuTxSJ
DhWRSrRasVznIcrWKmRfwtLwy5/4IeY+4BTlmdEGH3zishugzUV0+ApNhIx3hFMB
Vl7gX3Jt0iKEL5MKtOZRiV6FppGDVN9SIuDWQNymjfAZRp1IUuu69AemN2g4S5yF
A1Se2T2sJd1UId2h5bK/55UxHtitGfrgr3niuKH8L+D+KliqapNf0yWphgSVX6KD
bXTZckD8x0KOcMrXDOEqnkgyBiXmuQblfF9kiHXIyb3mdRWRfHG5VGHXBR21pUO8
Hg+0iK++kxVrCT8d9LNM+nbPQpMLUIEpVidQXkCsQ9sH1JS06BhHPlChArQ53jO6
N6wwHYAYh7FUii8WTKcFpOy5/BnNySIlnkYWvUJ5kq9GnPx6Q2twWnQSrWCpd0gh
1VD6j1PASRgHthzBqNzYBNOmTK79j1eZb0i6Udao4DmhF2OmZcMkGAYRK9oCZbT8
77NA26RZh3u2y9iaDfg+nIEsGYPMKcIfof5Sy42CZKdik4lp8a6AUKicJY4DQ3dK
sADWCjMX0LCXyFH5KO4Qnzqy40I/cgOJok+I0nrApYBLJCsqDTzCqJewG9CPFQiV
1raFSjWPcRC7Y1CRO7++oxJwDj96lzUYaoTv37cLueycQsXbV0XESMd3a8qLyNND
w2/xCLnnzDcLhb9XKT1b5TrlSDgi2MCfCurEuF2UjFdUMqdqqUmB8kVKrmzazTj5
cMcJjbJ7F1eFT5W6mqcI8cA1Jhtbc8M6Fe2z9er16wcQuOM4L0+tYkJrqx8OgsiT
wOuY0D2Hk2qS2PFDGdLqByDr3sE7BLWNfZ9hW8MDMi8QPvaNABedNm4Hi0tfYA+5
8KG7BjxOZNTPiI0kHC4kf3Ugy79Epx/3tMdrirKzRnmqArk8/acEKdJYws664XAR
WLAwAEFv7k/F4W5fTKyCuNho1VpSdKIDzvhHirnebuAytdcfAiFzhO/TeDkq76MB
vSB7I5QYwe4Nu0UaIoHWk0imu0JcnhQgFwSua1rf2jqKBAm7ByvP7jY6zLSP8jqq
thFxaZSak2y/sPB0J+clxEqnolaup2u3eLdB29Q7sygrNsc1YXFqKpAK6Zg0xaNT
zcdbe5TtDPcoq+hs53rYZnEYj0kt1CuoGQqUghI4UBUICjk3KD5ldBfqkU2l8QPf
h9SL2EVtDrsekjNglYOld6LVR9Mi7rrxEwAPiVbJpj2eYFUjDHGUXvG7rDUYYbjL
bZlt3rTOZlp/Q/zmGAfa4ASZbITutbMwE6DJe47jYzWo1oAQmnrJYEs7KaeqgzGT
5wBmFJehx+Zc9lXx9RQv+jewXK40U9nkLjMSjrJvYYtWMzNTlDBLaBqp/D4gQr1r
9LUFQYfX6nGNCImB5w2RSg==
`pragma protect end_protected
