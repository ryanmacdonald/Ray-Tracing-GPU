
module begin
  input clk, rst,

  input logic 

end
