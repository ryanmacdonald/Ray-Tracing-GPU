


module reflector(








endmodule: reflector
