/*
module send_shadow(
  
  input clk, rst,

  input scache_to_sendshadow_valid;
  input scache_to_sendshadow_t scache_to_sendshadow_data;
  output scache_to_sendshadow_stall;

  

  ) ;

endmodule*/
