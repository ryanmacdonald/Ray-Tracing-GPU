`default_nettype none

module frame_buffer_handler(
    // interface with pixel buffer
    output logic pb_re,
    input logic pb_empty,
    input pixel_buffer_entry_t pb_data,
    // sram interface
    output logic sram_oe_b,
    output logic sram_we_b,
    output logic sram_ce_b,
    output logic [19:0] sram_addr,
    inout wire [15:0] sram_io,
    output logic sram_ub_b, sram_lb_b,
    // vga interface
    output logic HS, VS,
    output logic VGA_clk,
    output logic VGA_blank,
    output logic [23:0] VGA_RGB,
    //
    input logic stripes_sel,
    input logic sq_sel,
    input logic[9:0] sq_row, sq_col,
    input logic clk, rst
);

    logic sram_re_b;
    assign sram_oe_b = sram_re_b;

    assign sram_ce_b = 1'b0;

    logic [19:0] writer_addr, reader_addr;
    logic [15:0] writer_data, reader_data;
    logic writer_ub, writer_lb;
    logic reader_ub, reader_lb;

    assign reader_data = sram_io;

    assign reader_ub = 1'b1;
    assign reader_lb = 1'b1;

    assign sram_io = (~sram_we_b) ? writer_data : 16'bz;
    assign sram_addr = (~sram_re_b) ? reader_addr : writer_addr;
    assign sram_lb_b = (~sram_re_b) ? ~reader_lb : ~writer_lb;
    assign sram_ub_b = (~sram_re_b) ? ~reader_ub : ~writer_ub;

    fbh_writer writer(.*);
    fbh_reader reader(.*);

endmodule: frame_buffer_handler

module fbh_writer(
    // pixel buffer
    output logic pb_re,
    input logic pb_empty,
    input pixel_buffer_entry_t pb_data,
    // SRAM
    output logic sram_we_b,
    output logic [19:0] writer_addr,
    output logic [15:0] writer_data,
    output logic writer_ub, writer_lb,
    //
    input logic sram_re_b, // from reader
    input logic clk, rst
);

    logic first_write, second_write;
    assign second_write = ~first_write;

    assign sram_we_b = ~(sram_re_b & ~pb_empty);
    assign pb_re = second_write & ~sram_we_b;

    color_t pb_pixel;
    pixel_buffer_entry_t pb_PID;
    logic [18:0] PID_addr0, PID_addr1;
    assign pb_pixel = pb_data.color;
    assign pb_PID = pb_data.pixelID.pixelID;

    assign PID_addr0 = pb_PID + (pb_PID >> 1'b1);
    assign PID_addr1 = PID_addr0+1'b1;

    // TODO: make sure these are not swapped incorrectly
    assign writer_ub = ~pb_PID[0] | second_write;
    assign writer_lb = pb_PID[0] | first_write;

    always_comb begin
        case({first_write,pb_PID[0]}) // TODO: get bit 0 of pixelID specifically
			// chronological order
            2'b10: writer_data = {pb_pixel.red, pb_pixel.green};
            2'b00: writer_data = {pb_pixel.blue,  8'b0};
            2'b11: writer_data = {8'b0,           pb_pixel.red};
            2'b01: writer_data = {pb_pixel.green, pb_pixel.blue};
        endcase
    end

    assign writer_addr = (first_write) ? {1'b0, PID_addr0} : {1'b0, PID_addr1}; // TODO: MSB should flip for double frame buffer

    ff_ar_en #(1,1'b1) first_write_ff(.q(first_write), .d(~first_write), .en(~sram_we_b), .clk, .rst);

endmodule: fbh_writer

module fbh_reader(
    // to VGA
    output logic HS, VS,
    output logic VGA_clk,
    output logic VGA_blank,
    output logic [23:0] VGA_RGB,
    // to/from SRAM
    output logic sram_re_b,
    output logic [19:0] reader_addr,
    input logic [15:0] reader_data,
    //
    input logic stripes_sel,
    input logic sq_sel,
    input logic[9:0] sq_row, sq_col,
    input logic clk, rst
);

    // vga controller
    logic display_done;
    logic [9:0] vga_row;
    logic [9:0] vga_col;
    logic clk_25M;
    logic clk_50M;
    assign clk_50M = clk;
    vga vc(.*);    

    // fbh_active
    logic row_on_screen;
    logic fbh_active, flip_active_on, flip_active_off;
    assign flip_active_on = (vga_col == 10'h3fe & row_on_screen);
    assign flip_active_off = (vga_col == 10'h27e);
    ff_ar_en #(1,1'b0) fbh_active_ff(.q(fbh_active), .d(flip_active_on), .en(flip_active_on | flip_active_off), .clk, .rst);

    range_check #(.W(10)) row_rc(
        .is_between(row_on_screen),
        .val(vga_row), .low(10'd0), .high(10'd479));

    logic [3:0] abc_sr_q;
    logic [15:0] a_q, b_q, c_q;
    logic a_en, b_en, c_en;
    logic [2:0] stripes_color, square_color;

    // address counter
    logic addr_cnt_inc, addr_cnt_clr;
    assign addr_cnt_inc = fbh_active & (a_en | b_en | c_en);
    assign addr_cnt_clr = (vga_row == 10'd0 && vga_col == 10'h3fd);
    counter #(20,20'd0) addr_counter(.cnt(reader_addr), .inc(addr_cnt_inc), .clr(addr_cnt_clr), .clk, .rst);

    shifter #(4,4'b100) abc_sr(.q(abc_sr_q), .d(abc_sr_q[0]), .en(fbh_active), .clr(addr_cnt_clr), .clk, .rst);

    // a, b, and c registers
    assign a_en = abc_sr_q[2];
    assign b_en = abc_sr_q[1];
    assign c_en = abc_sr_q[0];
    assign sram_re_b = ~((a_en | b_en | c_en) & fbh_active);

    ff_ar_en #(16,16'd0) a_reg(.q(a_q), .d(reader_data), .en(a_en), .clk, .rst); // first two bytes of first pixel
    ff_ar_en #(16,16'd0) b_reg(.q(b_q), .d(reader_data), .en(b_en), .clk, .rst); // third byte of first and first byte of second
    ff_ar_en #(16,16'd0) c_reg(.q(c_q), .d(reader_data), .en(c_en), .clk, .rst); // last two bytes of second pixel

    // pixel mux
    logic pixel_mux_sel;
    logic flip_pixel_mux_sel;
    assign flip_pixel_mux_sel = (a_en | c_en) & fbh_active;

    ff_ar_en #(1,1'b0) pixel_mux_sel_ff(.q(pixel_mux_sel), .d(~pixel_mux_sel), .en(flip_pixel_mux_sel), .clk, .rst);

    // pixel reg
    logic [23:0] pixel_reg_q, pixel_reg_d;
    assign pixel_reg_d = (pixel_mux_sel) ? {a_q, b_q[15:8]} : {b_q[7:0], c_q};
    ff_ar_en #(24,24'd0) pixel_reg(.q(pixel_reg_q), .d(pixel_reg_d), .en(flip_pixel_mux_sel), .clk, .rst);

    stripes stripes_inst(.vga_color(stripes_color), .vga_row, .vga_col);
    square   square_inst(.vga_color(square_color),.vga_row, .vga_col, .sq_row, .sq_col);

    // VGA output
    assign VGA_RGB = (stripes_sel) ? { stripes_color[2],7'b0, stripes_color[1],7'b0, stripes_color[0],7'b0} :
		     ( sq_sel ? { square_color[2],7'b0, square_color[1],7'b0, square_color[0],7'b0} : pixel_reg_q);

endmodule: fbh_reader
