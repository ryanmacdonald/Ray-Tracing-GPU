


module reflector();








endmodule: reflector
