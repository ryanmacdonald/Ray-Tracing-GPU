/* The Teal Rime Tray Racer! */
// Paul Kennedy   <pmkenned>
// Ross Daly      <rdaly>
// Ryan MacDonald <rmacdona>

module trtr();

endmodule
