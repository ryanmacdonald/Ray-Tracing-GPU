/* 
  Fully pipelined 1/1 intersection unit.
  Takes in a cacheline (Matrix + translate)
  A ray_vec
  and does a intersection test with them (t_int > epsilon && bari_test)  NO MAX test

*/

module int_unit(


  );


endmodule
